module VGA_Controller ();

endmodule // VGA_Controller
