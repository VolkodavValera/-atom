//`include "vga_avalon.svh"

module mem2vga (
	// Clock
	clk,

	// Asynchronous reset active low
	rst_n,

/*	// AVALON Interface
	address,
	read,
	readdata,
	write,
	writedata,
*/
	// SDRAM Interface
/*	sdram_addr,
	sdram_ba,
	sdram_cas_n,
	sdram_cke,
	sdram_cs_n,
	sdram_dq,
	sdram_dqm,
	sdram_ras_n,
	sdram_we_n,
	sdram_clk,
*/
	// VGA Interface
	VGA_HS,
	VGA_VS,
	VGA_R,
	VGA_G,
	VGA_B,

	// Other
	SW,
	LED,

	// arinc
	write,
	arinc_date,
	empty
);

/*------------------------------------------------------*/
/*						Parameters						*/
/*------------------------------------------------------*/
	parameter ADDRESS_WIDTH		= 3;
	localparam WAIT_ARINC		= 0;
	localparam FIFO_ARINC_FULL 	= 1;
	localparam READ_DATA		= 2;
	localparam FIFO_ARINC_EMPTY	= 3;


/*------------------------------------------------------*/
/*						Input							*/
/*------------------------------------------------------*/
	input							clk;
	input							rst_n;
/* 	input [ADDRESS_WIDTH - 1:0]		address;
	input							read;
	input							write;
	input [31:0]					writedata;
*/
	input [1:0]						SW;

	input 							write;
	input [31:0]					arinc_date;

/*------------------------------------------------------*/
/*						Output							*/
/*------------------------------------------------------*/
//	output 	[31:0]					readdata;
/*
    output	[12:0]					sdram_addr;
	output	[1:0]					sdram_ba;
	output							sdram_cas_n;
	output							sdram_cke;
	output							sdram_cs_n;
	output	[1:0]					sdram_dqm;
	output							sdram_ras_n;
	output							sdram_we_n;
	output							sdram_clk;
*/
	output							VGA_HS;					//	VGA H_SYNC
	output							VGA_VS;					//	VGA V_SYNC
	output	[3:0]					VGA_R;   				//	VGA Red[3:0]
	output	[3:0]					VGA_G;	 				//	VGA Green[3:0]
	output	[3:0]					VGA_B;   				//	VGA Blue[3:0]

	output 	[9:0]					LED;

	output 							empty;


/*------------------------------------------------------*/
/*						Inout							*/
/*------------------------------------------------------*/
//	inout	[15:0]					sdram_dq;

/*------------------------------------------------------*/
/*						Variables						*/
/*------------------------------------------------------*/

	// PLL signals
	// ---------------------------------------------------
	wire 							clk_sys;
	wire 							clk_vga;
	wire 	[1:0]					clk_pll;

	// FIFO A708
	// ---------------------------------------------------
	wire 							fifo_a708_empty;
	wire 							fifo_a708_full;
	wire 							fifo_a708_write;
	wire 							fifo_a708_read;
	wire 	[31:0]					fifo_a708_input_date;
	wire 	[31:0]					fifo_a708_output_date;

	logic 							package_arrived;
	logic 							package_arrived_ff;
	wire 							addr_gen_read;

	// FIFO NIOS II
	// ---------------------------------------------------
/*	wire 							fifo_nios_empty;
	wire 							fifo_nios_full;
	wire 							fifo_nios_write;
	wire 							fifo_nios_read;
	wire 	[31:0]					fifo_nios_input_date;
	wire 	[31:0]					fifo_nios_output_date;

	// FIFO VGA
	// ---------------------------------------------------
	wire 							fifo_vga_empty;
	wire 							fifo_vga_full;
	wire 							fifo_vga_write;
	wire 							fifo_vga_read;
	wire 	[2:0]					fifo_vga_input_date;
	wire 	[2:0]					fifo_vga_output_date;
*/
	// SDRAM Interface
	// ---------------------------------------------------
/*	wire 	[24:0]					sdram_write_address;
	wire 	[15:0]					sdram_write_data;
	wire 							sdram_write_enable;

	wire 	[24:0]					sdram_read_address;
	wire 	[15:0]					sdram_read_data;
	wire 							sdram_read_enable;
	wire 							sdram_read_ready;

	wire 							sdram_busy;
*/
	// RAM
	logic 	[2:0] 					RAM_Q;
	wire 	[18:0]					RAM_ADDR;
	wire 	[18:0]					ram_read_address;
	wire 	[18:0]					ram_write_address;
	wire 							ram_write;

	// ROM
	wire 	[11:0]					ROM_Q;
	wire 	[2:0]					ROM_ADDR;


	// Mashine
	logic	[2:0]					state;

	// Avalon
	wire 	[ADDRESS_WIDTH - 1:0]	address;
	wire							read;
	wire							write;
	wire 	[31:0]					writedata;
	wire 	[31:0]					readdata;

	logic 	[11:0] 					grad_gen_input;
	//logic 	[7:0]					angle;

/*------------------------------------------------------*/
/*						Сonnections						*/
/*------------------------------------------------------*/
	assign clk_sys = clk_pll[0];																	// System clock - 100 MHz
	assign sdram_clk = clk_pll[1];																	// Clock SDRAM - 100 MHZ + shift
	assign RAM_ADDR = ram_write ? ram_write_address : ram_read_address;								// If not write in RAM => read
	//assign ROM_ADDR = (RAM_Q);
	assign ROM_ADDR = (mem[ram_read_address]);

	assign fifo_a708_read = (package_arrived || package_arrived_ff || addr_gen_read) ? 1 : 0;		// If you received the entire package or read command from the module ADDR_GEN => Read FIFO
	assign fifo_a708_input_date = arinc_date;
	assign fifo_a708_write = write;
	assign empty = fifo_a708_empty;
	assign LED = (SW[0]) ? 10'h2AA : (SW[1]) ? 10'h1DD : 10'h3F1;

/*------------------------------------------------------*/
/*						Always blocks					*/
/*------------------------------------------------------*/

	// If FIFO=full => read header - 64 bits
	always_ff @(posedge clk_sys) begin
		if (fifo_a708_full) package_arrived <= 1'b1;
		else package_arrived <= 1'b0;

		package_arrived_ff <= package_arrived;
	end

	always_ff @(posedge clk_sys) begin
		if (!rst_n) grad_gen_input <= '0;
		else if (package_arrived_ff) grad_gen_input <= fifo_a708_output_date[31:20];
	end

	// RAM
	/*always_ff @ (posedge clk_sys) begin
		RAM_Q <= (mem[{ram_read_address}]);
	end*/


/*------------------------------------------------------*/
/*						Modules							*/
/*------------------------------------------------------*/
	/*SDRAM_Controller SDRAM (
			.wr_addr       (sdram_write_address),
			.wr_data       (sdram_write_data),
			.wr_enable     (sdram_write_enable),

			.rd_addr       (sdram_read_address),
			.rd_data       (sdram_read_data),
			.rd_ready      (sdram_read_ready),
			.rd_enable     (sdram_read_enable),

			.busy          (sdram_busy),
			.rst_n         (rst_n),
			.clk           (clk_sys),

			// SDRAM SIDE
			.addr          (sdram_addr),
			.bank_addr     (sdram_ba),
			.data          (sdram_dq),
			.clock_enable  (sdram_cke),
			.cs_n          (sdram_cs_n),
 			.ras_n         (sdram_ras_n),
			.cas_n         (sdram_cas_n),
			.we_n          (sdram_we_n),
			.data_mask_low (sdram_dqm[0]),
 			.data_mask_high(sdram_dqm[1]));*/

	VGA_Controller VGA (
			.clk_vga(clk_vga),
			.rst_n(rst_n),

			// Read date
			.address_vga(ram_read_address),
			.data(ROM_Q),

			// VGA SIDE
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.SW(SW));

	// Writing to RAM
	Generate_Addr ADDR_GEN (
		.clk(clk_sys),
		.rst_n(rst_n),
		.angle(grad_gen_input),
		.ADDR_RAM_WRITE(ram_write_address),
		.RAM_WRITE(ram_write),
		.FIFO_READ(addr_gen_read));
/*
	// Converting relative angle to absolute from 0 to 180
	Floating_point Grad_Gen (
		.clk(clk_sys),
		.rst_n(rst_n),
		.in_arinc(grad_gen_input),
		.graf_angle(angle));
*/
/*------------------------------------------------------*/
/*						RAM								*/
/*------------------------------------------------------*/
	/*altsyncram	RAM_DISPLEY (
				.address_a (RAM_ADDR),
				.clock0 (clk_sys),
				.data_a (fifo_a708_output_date),
				.wren_a (ram_write),
				.q_a (RAM_Q),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.address_b (1'b1),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_b (1'b1),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_b (1'b0));
	defparam
		RAM_DISPLEY.clock_enable_input_a = "BYPASS",
		RAM_DISPLEY.clock_enable_output_a = "BYPASS",
		RAM_DISPLEY.intended_device_family = "MAX 10",
		RAM_DISPLEY.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
		RAM_DISPLEY.lpm_type = "altsyncram",
		RAM_DISPLEY.numwords_a = 307200,
		RAM_DISPLEY.operation_mode = "SINGLE_PORT",
		RAM_DISPLEY.outdata_aclr_a = "NONE",
		RAM_DISPLEY.outdata_reg_a = "CLOCK0",
		RAM_DISPLEY.power_up_uninitialized = "FALSE",
		RAM_DISPLEY.read_during_write_mode_port_a = "NEW_DATA_NO_NBE_READ",
		RAM_DISPLEY.widthad_a = 19,
		RAM_DISPLEY.width_a = 3,
		RAM_DISPLEY.width_byteena_a = 1;
*/

/*------------------------------------------------------*/
/*						FIFO							*/
/*------------------------------------------------------*/

	// write ARINC708 -> read NIOS II 						- 1600 bits = 50 * 32 bits
	dcfifo	fifo_a708 (
			.aclr (~rst_n),
			.data (fifo_a708_input_date),
			.rdclk (clk_sys),
			.rdreq (fifo_a708_read),
			.wrclk (clk),
			.wrreq (fifo_a708_write),
			.q (fifo_a708_output_date),
			.rdempty (fifo_a708_empty),
			.wrfull (fifo_a708_full)
			);

	defparam
			fifo_a708.intended_device_family = "MAX 10",
			fifo_a708.lpm_numwords = 50,
			fifo_a708.lpm_showahead = "OFF",
			fifo_a708.lpm_type = "dcfifo",
			fifo_a708.lpm_width = 32,
			fifo_a708.lpm_widthu = 6,
			fifo_a708.overflow_checking = "ON",
			fifo_a708.rdsync_delaypipe = 4,
			fifo_a708.read_aclr_synch = "OFF",
			fifo_a708.underflow_checking = "ON",
			fifo_a708.use_eab = "ON",
			fifo_a708.write_aclr_synch = "OFF",
			fifo_a708.wrsync_delaypipe = 4;


	// write NIOS II -> read SDRAM Controller 				- 1 row - 640 * 3 bits = 60 * 32 bits
/*	scfifo fifo_nios
		(
			.rdreq(fifo_nios_read),
			.aclr(~rst_n),
			.sclr(),
			.clock(clk_sys),
			.wrreq(fifo_nios_write),
			.data(fifo_nios_input_date),
			.usedw(),
			.empty(fifo_nios_empty),
			.full(fifo_nios_full),
			.q(fifo_nios_output_date)
		);

	defparam
			fifo_nios.add_ram_output_register = "OFF",
			fifo_nios.intended_device_family = "MAX 10",
			fifo_nios.lpm_numwords = 60,
			fifo_nios.lpm_showahead = "OFF",
			fifo_nios.lpm_type = "scfifo",
			fifo_nios.lpm_width = 32,
			fifo_nios.lpm_widthu = 6,
			fifo_nios.overflow_checking = "ON",
			fifo_nios.underflow_checking = "ON";

*/
	// write SDRAM Controller -> read VGA Controller 		- 1 row - 640 * 3 bits
/*	dcfifo	fifo_vga (
			.aclr (~rst_n),
			.data (fifo_vga_input_date),
			.rdclk (clk_vga),
			.rdreq (fifo_vga_read),
			.wrclk (clk_sys),
			.wrreq (fifo_vga_write),
			.q (fifo_vga_output_date),
			.rdempty (fifo_vga_empty),
			.wrfull (fifo_vga_full)
			);

	defparam
			fifo_vga.intended_device_family = "MAX 10",
			fifo_vga.lpm_numwords = 640,
			fifo_vga.lpm_showahead = "OFF",
			fifo_vga.lpm_type = "dcfifo",
			fifo_vga.lpm_width = 3,
			fifo_vga.lpm_widthu = 6,
			fifo_vga.overflow_checking = "ON",
			fifo_vga.rdsync_delaypipe = 4,
			fifo_vga.read_aclr_synch = "OFF",
			fifo_vga.underflow_checking = "ON",
			fifo_vga.use_eab = "ON",
			fifo_vga.write_aclr_synch = "OFF",
			fifo_vga.wrsync_delaypipe = 4;

*/
/*------------------------------------------------------*/
/*						PLL								*/
/*------------------------------------------------------*/
	altpll	PLL_VGA (
				.inclk (clk),
				.clk (clk_vga),
				.areset (1'b0),
				.clkena ({6{1'b1}}),
				.clkswitch (1'b0),
				.configupdate (1'b0),
				.extclkena ({4{1'b1}}),
				.fbin (1'b1),
				.pfdena (1'b1),
				.phasecounterselect ({4{1'b1}}),
				.phasestep (1'b1),
				.phaseupdown (1'b1),
				.pllena (1'b1),
				.scanaclr (1'b0),
				.scanclk (1'b0),
				.scanclkena (1'b1),
				.scandata (1'b0),
				.scanread (1'b0),
				.scanwrite (1'b0));
	defparam
		PLL_VGA.bandwidth_type = "AUTO",
		PLL_VGA.clk0_divide_by = 2000,
		PLL_VGA.clk0_duty_cycle = 50,
		PLL_VGA.clk0_multiply_by = 1007,
		PLL_VGA.clk0_phase_shift = "0",
		PLL_VGA.compensate_clock = "CLK0",
		PLL_VGA.inclk0_input_frequency = 20000,
		PLL_VGA.intended_device_family = "MAX 10",
		PLL_VGA.lpm_type = "altpll",
		PLL_VGA.operation_mode = "NORMAL",
		PLL_VGA.pll_type = "AUTO",
		PLL_VGA.port_clk0 = "PORT_USED",
		PLL_VGA.width_clock = 1;


	altpll	PLL_SDRAM (
				.inclk (clk),
				.clk (clk_pll),
				.areset (1'b0),
				.clkena ({6{1'b1}}),
				.clkswitch (1'b0),
				.configupdate (1'b0),
				.extclkena ({4{1'b1}}),
				.fbin (1'b1),
				.pfdena (1'b1),
				.phasecounterselect ({4{1'b1}}),
				.phasestep (1'b1),
				.phaseupdown (1'b1),
				.pllena (1'b1),
				.scanaclr (1'b0),
				.scanclk (1'b0),
				.scanclkena (1'b1),
				.scandata (1'b0),
				.scanread (1'b0),
				.scanwrite (1'b0));
	defparam
		PLL_SDRAM.bandwidth_type = "AUTO",
		PLL_SDRAM.clk0_divide_by = 36,
		PLL_SDRAM.clk0_duty_cycle = 50,
		PLL_SDRAM.clk0_multiply_by = 103,
		PLL_SDRAM.clk0_phase_shift = "0",
		PLL_SDRAM.clk1_divide_by = 36,
		PLL_SDRAM.clk1_duty_cycle = 50,
		PLL_SDRAM.clk1_multiply_by = 103,
		PLL_SDRAM.clk1_phase_shift = "-3000",
		PLL_SDRAM.compensate_clock = "CLK0",
		PLL_SDRAM.inclk0_input_frequency = 20000,
		PLL_SDRAM.intended_device_family = "MAX 10",
		PLL_SDRAM.lpm_type = "altpll",
		PLL_SDRAM.operation_mode = "NORMAL",
		PLL_SDRAM.pll_type = "AUTO",
		PLL_SDRAM.port_clk0 = "PORT_USED",
		PLL_SDRAM.port_clk1 = "PORT_USED",
		PLL_SDRAM.width_clock = 2;

/*------------------------------------------------------*/
/*						ROM								*/
/*------------------------------------------------------*/
	altsyncram	ROM_Palitra (
				.address_a (ROM_ADDR),
				.clock0 (clk_sys),
				.q_a (ROM_Q),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.address_b (1'b1),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_a ({12{1'b1}}),
				.data_b (1'b1),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_a (1'b0),
				.wren_b (1'b0));
	defparam
		ROM_Palitra.address_aclr_a = "NONE",
		ROM_Palitra.clock_enable_input_a = "BYPASS",
		ROM_Palitra.clock_enable_output_a = "BYPASS",
		ROM_Palitra.init_file = "./source/palitra.hex",
		ROM_Palitra.intended_device_family = "MAX 10",
		ROM_Palitra.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
		ROM_Palitra.lpm_type = "altsyncram",
		ROM_Palitra.numwords_a = 8,
		ROM_Palitra.operation_mode = "ROM",
		ROM_Palitra.outdata_aclr_a = "NONE",
		ROM_Palitra.outdata_reg_a = "CLOCK0",
		ROM_Palitra.widthad_a = 3,
		ROM_Palitra.width_a = 12,
		ROM_Palitra.width_byteena_a = 1;

logic [2:0] mem [30720] =
	'{
		3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b111, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b001, 3'b110, 3'b001, 3'b101, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b101, 3'b011, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b001,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b000,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b001, 3'b111, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b000,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b001, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b000, 3'b010, 3'b101, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b111, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b111, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b011, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b000, 3'b100,
		3'b000, 3'b000, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b111,
		3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000,
		3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b110, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b001, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b001, 3'b001, 3'b111, 3'b000, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b110, 3'b000, 3'b010, 3'b000,
		3'b001, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011,
		3'b101, 3'b110, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011, 3'b000,
		3'b000, 3'b011, 3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b010, 3'b000, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b111, 3'b111, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b011, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b000, 3'b101, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b000, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b111, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b111, 3'b001, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111,
		3'b000, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b101, 3'b110, 3'b101,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b001, 3'b110, 3'b000, 3'b000,
		3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b111, 3'b110, 3'b010, 3'b001, 3'b011, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b011, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b000, 3'b011, 3'b001, 3'b010, 3'b000, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b000, 3'b001, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b000, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b110, 3'b101, 3'b111,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b001, 3'b110, 3'b110, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111,
		3'b111, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b000, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b110, 3'b101, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b111, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b011,
		3'b000, 3'b010, 3'b110, 3'b101, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b000, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b011, 3'b110, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b101, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b000, 3'b001, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b001, 3'b111, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110,
		3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000,
		3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b101, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101,
		3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b110, 3'b010, 3'b101, 3'b101, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b001, 3'b001, 3'b111, 3'b001,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b101, 3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b101, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b000, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b101, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b111, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b011, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b000, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b111,
		3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000, 3'b111, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101,
		3'b100, 3'b101, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b111, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b111,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b110, 3'b011, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b011, 3'b101, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b110, 3'b001, 3'b111, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b101, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b110, 3'b110, 3'b110, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b001, 3'b101, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b001, 3'b001, 3'b101, 3'b100, 3'b110, 3'b011, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b000, 3'b110, 3'b100, 3'b111, 3'b110, 3'b111, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b000, 3'b000, 3'b001, 3'b101, 3'b010, 3'b101, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b001, 3'b000, 3'b000, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b011, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b000, 3'b000, 3'b100, 3'b101, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b001, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b011, 3'b010, 3'b000, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b011, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b001, 3'b101, 3'b111, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b011, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b111, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b111, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b111, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b011, 3'b101, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b011, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b101, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b111, 3'b101, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b111, 3'b111, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b111, 3'b100, 3'b111, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b101, 3'b100, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b110, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b010, 3'b110, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b000,
		3'b000, 3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b111, 3'b111, 3'b010, 3'b111, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b011, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b001, 3'b000, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b101, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b010, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b001, 3'b000, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b101, 3'b011, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b000, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b010, 3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b111, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b001, 3'b001, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b110, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b011, 3'b000,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b011, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b101, 3'b111, 3'b000, 3'b010, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b111, 3'b000, 3'b010,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b111, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b000, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b101, 3'b101, 3'b010, 3'b001, 3'b011, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b111, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b001, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b000, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b011, 3'b000, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b000, 3'b101, 3'b101, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b111, 3'b001, 3'b010, 3'b100, 3'b001, 3'b101, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b101, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b011, 3'b011, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b000, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b011, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b000, 3'b101, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b011, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b000, 3'b100, 3'b000, 3'b110, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000, 3'b111, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b101, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b011, 3'b101, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b011, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b011, 3'b000, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b101, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b101, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b010, 3'b000, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b111, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b001, 3'b000, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001, 3'b111,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b111, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b001, 3'b111, 3'b111, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b110, 3'b011, 3'b101, 3'b011, 3'b100, 3'b001, 3'b011, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b000, 3'b111, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b101, 3'b101, 3'b001, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b111,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b101, 3'b010, 3'b011, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b101, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b000, 3'b110, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b111, 3'b010, 3'b100, 3'b011, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111,
		3'b010, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b100, 3'b111, 3'b011, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b101, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b000, 3'b001, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b000, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b011, 3'b000, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b101,
		3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b011,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b000, 3'b001, 3'b100, 3'b110, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b011, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b010, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b101, 3'b101, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b101, 3'b110, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b111, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b111, 3'b010, 3'b100, 3'b001, 3'b101, 3'b110, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100,
		3'b000, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b011, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111,
		3'b111, 3'b000, 3'b000, 3'b100, 3'b011, 3'b000, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b000, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b011, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b001,
		3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b011, 3'b111, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b111, 3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b010, 3'b000, 3'b110, 3'b011, 3'b011, 3'b000, 3'b111, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b111, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011,
		3'b011, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b001, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000, 3'b101, 3'b101, 3'b000, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b100, 3'b111, 3'b101, 3'b101, 3'b000, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110,
		3'b011, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b000, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b001,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b001, 3'b001, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b101, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101,
		3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b000, 3'b010, 3'b001, 3'b110, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b111, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b000, 3'b010, 3'b001, 3'b101, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b001, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b011, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100
	};


endmodule: mem2vga
