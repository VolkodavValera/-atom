logic [2:0] mem [307200] =
	'{
		3'b001, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b111, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011,
		3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b111,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b101, 3'b010, 3'b010, 3'b001, 3'b000, 3'b111, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b111, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110,
		3'b110, 3'b100, 3'b000, 3'b101, 3'b111, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b001, 3'b000, 3'b010, 3'b000,
		3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b001, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b010,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b111, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001,
		3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b001, 3'b001, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b000, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b110, 3'b010, 3'b011, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b101, 3'b110, 3'b010, 3'b011, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b111, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b011,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b010, 3'b011, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b110, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b110, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b011, 3'b100, 3'b110, 3'b010,
		3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b000, 3'b101, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b111, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b111, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b000, 3'b101, 3'b001, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b110, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b111, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b000, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b111, 3'b111, 3'b111, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b001, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111,
		3'b111, 3'b000, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b110, 3'b110, 3'b001, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b000, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b010, 3'b010, 3'b111,
		3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b101, 3'b010, 3'b101, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b111, 3'b101, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b110, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b101, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b011, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100,
		3'b011, 3'b100, 3'b011, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b101, 3'b011, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b111, 3'b110, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b111, 3'b110, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b110, 3'b011, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b111, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b011, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110,
		3'b100, 3'b101, 3'b111, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b001, 3'b011, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101, 3'b010, 3'b111, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100,
		3'b010, 3'b101, 3'b000, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b111, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b111, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010,
		3'b000, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b111, 3'b111, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b001, 3'b011, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b101, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b011, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b011, 3'b001, 3'b001, 3'b011, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b101, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b010, 3'b011, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b110, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b101, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b001, 3'b011, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b011, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b110, 3'b000, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b000, 3'b110, 3'b011, 3'b010, 3'b011, 3'b111, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b110, 3'b101, 3'b001, 3'b101, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b010, 3'b001, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110,
		3'b111, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b000, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b111, 3'b101, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b001, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b011, 3'b110, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b101, 3'b001, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b111, 3'b001, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b011, 3'b010, 3'b110, 3'b011, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111,
		3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b011, 3'b110, 3'b110, 3'b110, 3'b000, 3'b011, 3'b111, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b111, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b000, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b011, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100,
		3'b011, 3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111,
		3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b011,
		3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b000, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101,
		3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b111, 3'b011, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b101, 3'b001, 3'b110, 3'b100, 3'b011, 3'b001, 3'b001, 3'b110, 3'b100,
		3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b111, 3'b001, 3'b010, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b110, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b001, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b101, 3'b010, 3'b101, 3'b000, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b101, 3'b000, 3'b011, 3'b100, 3'b110, 3'b101, 3'b000, 3'b001, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b110, 3'b001, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b101, 3'b001,
		3'b111, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b111, 3'b011, 3'b100, 3'b111, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b001, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b101, 3'b011, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b011, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b001,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000, 3'b111, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b101, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b111, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b101, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b010, 3'b101, 3'b010,
		3'b110, 3'b110, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b000, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b111,
		3'b000, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b011, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b101, 3'b001,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b011,
		3'b101, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b001, 3'b101, 3'b110, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b001, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b010, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b000, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b001,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b011, 3'b000, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b001, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b111, 3'b101, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b111, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b011, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b101, 3'b101, 3'b111, 3'b100, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b110, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b011, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b110, 3'b101, 3'b010,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b110, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b000, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b001,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b000, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111,
		3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b000, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b001, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b011, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001,
		3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b101, 3'b100, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b011, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b110, 3'b111, 3'b000, 3'b010, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111,
		3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b011, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b011,
		3'b000, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011, 3'b010, 3'b001, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b000, 3'b011, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b011, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b110, 3'b010, 3'b011,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b001, 3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b011, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b111, 3'b000, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b111, 3'b110, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b101, 3'b011, 3'b101, 3'b000, 3'b001, 3'b101, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b001, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b001, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b010, 3'b010, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b101,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b000, 3'b001, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010,
		3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b101, 3'b011, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b101, 3'b010, 3'b101, 3'b101, 3'b100, 3'b011, 3'b001, 3'b010, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010,
		3'b011, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b001, 3'b011, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b001, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b101, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b001, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b011,
		3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b011, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111,
		3'b011, 3'b110, 3'b010, 3'b011, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b001, 3'b110, 3'b110, 3'b101, 3'b100, 3'b101, 3'b101, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b111, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b011, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b000, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b101, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b110, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b101, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b001, 3'b001, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b111, 3'b000, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b101, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b000, 3'b101, 3'b011, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b000, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b011, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b101, 3'b010, 3'b111, 3'b010, 3'b001, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b001, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b111, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b000, 3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010,
		3'b010, 3'b110, 3'b111, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b011, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b011, 3'b011, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b000, 3'b001,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b000, 3'b011, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b011, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b001, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b000, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b000, 3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b101, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b000, 3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b111, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b000, 3'b011, 3'b100, 3'b101, 3'b010, 3'b001, 3'b110, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b111, 3'b100, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110,
		3'b110, 3'b111, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b110, 3'b000, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b101,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b111, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b001, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b011, 3'b000, 3'b010, 3'b110,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b101, 3'b001, 3'b101, 3'b000, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b111,
		3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b011, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b000, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b011, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b111, 3'b001, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b101, 3'b101, 3'b111, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b011, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b111, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b001, 3'b101, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b101, 3'b010, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110,
		3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b111, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b001, 3'b101, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b010, 3'b101, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b000, 3'b110, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b110, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b001, 3'b010,
		3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b011, 3'b110, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111, 3'b110, 3'b101, 3'b110, 3'b010, 3'b101,
		3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b111, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 3'b110, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b000, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b000, 3'b011, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b000, 3'b110, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b011, 3'b001, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b011, 3'b011, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b000, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b001, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b001, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b101, 3'b000, 3'b111, 3'b010,
		3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b001,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b111, 3'b010, 3'b101, 3'b010, 3'b001,
		3'b000, 3'b001, 3'b110, 3'b000, 3'b100, 3'b111, 3'b000, 3'b010, 3'b110, 3'b011, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b000, 3'b110,
		3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b011, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b001, 3'b101, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b011, 3'b010, 3'b100, 3'b000, 3'b011, 3'b110, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b011, 3'b011, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b001,
		3'b011, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b000,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b001, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b000, 3'b010, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b000, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b000, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b111, 3'b111, 3'b110, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b011, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b000, 3'b101, 3'b011, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010,
		3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b110, 3'b111, 3'b101, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b011, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b010, 3'b111, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b001, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b110, 3'b101,
		3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b110, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b011, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000, 3'b101, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010,
		3'b111, 3'b011, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b110, 3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b001, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b001, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b011,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b101, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b010, 3'b001, 3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b010, 3'b011, 3'b110, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b010, 3'b110, 3'b110, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b000, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b111, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b111, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b011, 3'b110, 3'b101, 3'b100, 3'b101, 3'b001, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b000, 3'b010,
		3'b111, 3'b001, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100,
		3'b111, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b001, 3'b000, 3'b110, 3'b101, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b011, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b000, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b011, 3'b111, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b110, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b101, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b101, 3'b010,
		3'b110, 3'b101, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b100, 3'b011, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b111, 3'b100, 3'b101, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b110, 3'b000, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b110, 3'b110, 3'b110,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b111, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b011, 3'b100, 3'b101, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b101, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b011, 3'b001, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b111, 3'b101, 3'b100, 3'b010,
		3'b000, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b001, 3'b001, 3'b000, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b001, 3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b000, 3'b101, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b000, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b111, 3'b111, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b000, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b001, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b001, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b011, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111,
		3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b110, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b000, 3'b110, 3'b011, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b111, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b001, 3'b110,
		3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b001, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b001, 3'b111, 3'b111,
		3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b011, 3'b001, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b101, 3'b000, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b011, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b001, 3'b000, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b001, 3'b101, 3'b000, 3'b110, 3'b011, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b111, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b101, 3'b110, 3'b010, 3'b110, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b101, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b000, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b111, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b111, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b101, 3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b000, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b010, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b001, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b110, 3'b010, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b011, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b111, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b111, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b111, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b101, 3'b011, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b111, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b111, 3'b111, 3'b110, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b011, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b101, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b110, 3'b101, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b111, 3'b100, 3'b010, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b101, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b111, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b111, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b010, 3'b111, 3'b000, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b001, 3'b010,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b001, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b111, 3'b110, 3'b110, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b011,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b101, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b001, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b001, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b111, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b011, 3'b010,
		3'b111, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b011,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b101, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b101, 3'b101, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b111, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b011,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b111, 3'b001, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010,
		3'b101, 3'b111, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b001, 3'b010, 3'b000, 3'b111, 3'b010, 3'b011, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b111, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101,
		3'b000, 3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b011, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b001, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b101, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b111, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b011,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b010, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b000, 3'b101, 3'b000, 3'b111, 3'b100, 3'b101, 3'b111, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b010, 3'b000, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b011,
		3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b110, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b101, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101,
		3'b110, 3'b011, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b001, 3'b110, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b101, 3'b011, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b110, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b011, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b111, 3'b001,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b000, 3'b111, 3'b101, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b011, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011,
		3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b111, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b011,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b011, 3'b001, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b101, 3'b111, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b001, 3'b101, 3'b001, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010,
		3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b011, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b011, 3'b011, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b111, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b000, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b101, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b011, 3'b011, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b111, 3'b111, 3'b110, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b000, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b000, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010,
		3'b101, 3'b010, 3'b001, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b110, 3'b101, 3'b000, 3'b101, 3'b110, 3'b111, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b010, 3'b111, 3'b011, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b001, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b000, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100,
		3'b010, 3'b101, 3'b000, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001, 3'b000, 3'b000, 3'b101, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b001, 3'b110, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b001, 3'b110, 3'b110, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b110, 3'b000, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b111, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b101, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b000,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b101, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b000, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b000, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b011, 3'b000, 3'b101, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b101, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b001, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b110, 3'b101, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b101, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b101, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b101, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b000, 3'b111, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111,
		3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b001, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b101,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b011, 3'b010, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110,
		3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b011, 3'b011, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b000, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b111, 3'b101, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b011, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b011, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b101, 3'b101, 3'b111, 3'b010,
		3'b010, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011,
		3'b010, 3'b100, 3'b000, 3'b110, 3'b111, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b110, 3'b000, 3'b001,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b010,
		3'b001, 3'b011, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b011, 3'b011, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b010, 3'b110, 3'b110, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b000, 3'b101, 3'b010, 3'b000, 3'b110,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b101, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b111, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b011, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b101, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b011, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b110, 3'b000, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b000, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b011, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110,
		3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b101,
		3'b010, 3'b000, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b101,
		3'b010, 3'b011, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b001, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b011, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b111, 3'b010,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b110, 3'b001, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b101, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b101, 3'b001, 3'b101, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b110, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b111, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b001,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b111, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b011,
		3'b010, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b101, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b001, 3'b011, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b111, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b101, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b111, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b010, 3'b101, 3'b000, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b001, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000, 3'b111, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b001,
		3'b001, 3'b110, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b011, 3'b000, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b001, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b000,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b001, 3'b011, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b000, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b001, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b111, 3'b001, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b111, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000,
		3'b001, 3'b001, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b001, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b001, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100,
		3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b111, 3'b101, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001, 3'b000, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b101, 3'b011, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b011, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b101, 3'b011, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b011, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b001, 3'b011, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b000, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b111, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b101, 3'b100, 3'b000, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b010, 3'b011, 3'b111, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b110, 3'b000, 3'b000, 3'b001, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b000, 3'b011, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b011,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b000, 3'b000, 3'b110, 3'b101, 3'b101,
		3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b111, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b011, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b011, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011, 3'b010, 3'b001, 3'b000, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b111, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b011, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b011, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b010, 3'b001, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b001, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b110, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100,
		3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b101, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b000, 3'b000, 3'b010, 3'b001, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b001, 3'b001, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b111, 3'b011, 3'b100, 3'b011, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b101, 3'b101, 3'b100, 3'b101, 3'b011, 3'b111, 3'b111, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b101, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b111,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b110,
		3'b010, 3'b000, 3'b010, 3'b000, 3'b110, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b001, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b101, 3'b000, 3'b001, 3'b001, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b101, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b011, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b111,
		3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b111, 3'b011, 3'b110, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b110, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b110, 3'b111, 3'b110, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b111, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b011, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011,
		3'b100, 3'b011, 3'b111, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b111, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b001, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b111, 3'b000, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111,
		3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b000, 3'b010, 3'b000, 3'b101, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b110, 3'b000,
		3'b000, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b000, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b111, 3'b110, 3'b001, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010, 3'b000, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b000, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b011, 3'b001, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b101, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b001, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101,
		3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b110, 3'b011, 3'b101, 3'b001, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b110, 3'b101,
		3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b111, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b001, 3'b000, 3'b111, 3'b000, 3'b010, 3'b010, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b000, 3'b000, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b011, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b111, 3'b001, 3'b010, 3'b111, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b001, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b101, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b000,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100,
		3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b110, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b011, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b011, 3'b011, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b101, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b011, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b110, 3'b110, 3'b010, 3'b110, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b000, 3'b001, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b110, 3'b111, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b111, 3'b110, 3'b000, 3'b111, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b011, 3'b010,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b011, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b111, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b001, 3'b110, 3'b001, 3'b101, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b101, 3'b011, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b001,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b000,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b001, 3'b111, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b000,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b001, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b000, 3'b010, 3'b101, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b111, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b111, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b011, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b000, 3'b100,
		3'b000, 3'b000, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b111,
		3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000,
		3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b110, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b001, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b001, 3'b001, 3'b111, 3'b000, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b110, 3'b000, 3'b010, 3'b000,
		3'b001, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011,
		3'b101, 3'b110, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011, 3'b000,
		3'b000, 3'b011, 3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b010, 3'b000, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b111, 3'b111, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b011, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b000, 3'b101, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b000, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b111, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b111, 3'b001, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111,
		3'b000, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b101, 3'b110, 3'b101,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b001, 3'b110, 3'b000, 3'b000,
		3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b111, 3'b110, 3'b010, 3'b001, 3'b011, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b011, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b000, 3'b011, 3'b001, 3'b010, 3'b000, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b000, 3'b001, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b000, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b110, 3'b101, 3'b111,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b001, 3'b110, 3'b110, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111,
		3'b111, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b000, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b110, 3'b101, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b111, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b011,
		3'b000, 3'b010, 3'b110, 3'b101, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b000, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b011, 3'b110, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b101, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b000, 3'b001, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b001, 3'b111, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110,
		3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000,
		3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b101, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101,
		3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b110, 3'b010, 3'b101, 3'b101, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b001, 3'b001, 3'b111, 3'b001,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b101, 3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b101, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b000, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b101, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b111, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b011, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b000, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b111,
		3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000, 3'b111, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101,
		3'b100, 3'b101, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b111, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b111,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b110, 3'b011, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b011, 3'b101, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b110, 3'b001, 3'b111, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b101, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b110, 3'b110, 3'b110, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b001, 3'b101, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b001, 3'b001, 3'b101, 3'b100, 3'b110, 3'b011, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b000, 3'b110, 3'b100, 3'b111, 3'b110, 3'b111, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b000, 3'b000, 3'b001, 3'b101, 3'b010, 3'b101, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b001, 3'b000, 3'b000, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b011, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b000, 3'b000, 3'b100, 3'b101, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b001, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b011, 3'b010, 3'b000, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b011, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b001, 3'b101, 3'b111, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b011, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b111, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b111, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b111, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b011, 3'b101, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b011, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b101, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b111, 3'b101, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b111, 3'b111, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b111, 3'b100, 3'b111, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b101, 3'b100, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b110, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b010, 3'b110, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b000,
		3'b000, 3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b111, 3'b111, 3'b010, 3'b111, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b011, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b001, 3'b000, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b101, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b010, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b001, 3'b000, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b101, 3'b011, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b000, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b010, 3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b111, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b001, 3'b001, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b110, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b011, 3'b000,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b011, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b101, 3'b111, 3'b000, 3'b010, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b111, 3'b000, 3'b010,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b111, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b000, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b101, 3'b101, 3'b010, 3'b001, 3'b011, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b111, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b001, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b000, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b011, 3'b000, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b000, 3'b101, 3'b101, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b111, 3'b001, 3'b010, 3'b100, 3'b001, 3'b101, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b101, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b011, 3'b011, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b000, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b011, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b000, 3'b101, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b011, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b000, 3'b100, 3'b000, 3'b110, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000, 3'b111, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b101, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b011, 3'b101, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b011, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b011, 3'b000, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b101, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b101, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b010, 3'b000, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b111, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b001, 3'b000, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001, 3'b111,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b111, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b001, 3'b111, 3'b111, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b110, 3'b011, 3'b101, 3'b011, 3'b100, 3'b001, 3'b011, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b000, 3'b111, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b101, 3'b101, 3'b001, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b111,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b101, 3'b010, 3'b011, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b101, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b000, 3'b110, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b111, 3'b010, 3'b100, 3'b011, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111,
		3'b010, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b100, 3'b111, 3'b011, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b101, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b000, 3'b001, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b000, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b011, 3'b000, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b101,
		3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b011,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b000, 3'b001, 3'b100, 3'b110, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b011, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b010, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b101, 3'b101, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b101, 3'b110, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b111, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b111, 3'b010, 3'b100, 3'b001, 3'b101, 3'b110, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100,
		3'b000, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b011, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111,
		3'b111, 3'b000, 3'b000, 3'b100, 3'b011, 3'b000, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b000, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b011, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b001,
		3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b011, 3'b111, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b111, 3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b010, 3'b000, 3'b110, 3'b011, 3'b011, 3'b000, 3'b111, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b111, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011,
		3'b011, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b001, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000, 3'b101, 3'b101, 3'b000, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b100, 3'b111, 3'b101, 3'b101, 3'b000, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110,
		3'b011, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b000, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b001,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b001, 3'b001, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b101, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101,
		3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b000, 3'b010, 3'b001, 3'b110, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b111, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b000, 3'b010, 3'b001, 3'b101, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b001, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b011, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b101,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b001, 3'b000, 3'b010, 3'b010,
		3'b001, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b111,
		3'b110, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b101, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b110, 3'b111, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b111, 3'b001, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b101, 3'b010, 3'b011, 3'b001, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b111, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b000, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b011, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b101, 3'b110, 3'b001, 3'b001,
		3'b010, 3'b000, 3'b111, 3'b111, 3'b010, 3'b110, 3'b000, 3'b100, 3'b011, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b011, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b011, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b101, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b111, 3'b011, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b101, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b011, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b011, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b011, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111,
		3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011, 3'b111, 3'b101,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b000, 3'b001, 3'b100, 3'b111,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b101, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b111,
		3'b001, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b111, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b011, 3'b110,
		3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b110, 3'b001, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b011, 3'b111, 3'b110, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b111, 3'b010, 3'b010, 3'b000, 3'b110, 3'b011, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b010,
		3'b001, 3'b000, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b000, 3'b101, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b001, 3'b010, 3'b101, 3'b001, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b111, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b011, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b000, 3'b110, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b001, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b001, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b111, 3'b100, 3'b010, 3'b000, 3'b111, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b101, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b110, 3'b001, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b111, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b000, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b101, 3'b011, 3'b101,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b011, 3'b110, 3'b101, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b000, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b100, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b001, 3'b000, 3'b111, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b110, 3'b011, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000,
		3'b001, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b111, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b101, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b101, 3'b010, 3'b000, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 3'b101, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b000, 3'b111, 3'b111, 3'b110, 3'b111,
		3'b011, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b111, 3'b000, 3'b001, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b000, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b101, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000,
		3'b000, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b011, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b000,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b001, 3'b000, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b011, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b000, 3'b111, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b001, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b110, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b001, 3'b001, 3'b001, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b111, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b001, 3'b000, 3'b101, 3'b010, 3'b010, 3'b110,
		3'b000, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b101, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b000, 3'b111, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b101, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b011, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b000, 3'b000, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b101, 3'b100, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b101, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010,
		3'b101, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b101, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b110, 3'b111, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b111, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b000, 3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b101, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b101, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b111,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b000, 3'b101, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b101,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b001, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b110, 3'b110, 3'b000,
		3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b101,
		3'b111, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b101, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b000, 3'b001, 3'b110, 3'b010, 3'b111, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b110, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b111, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b111,
		3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b011, 3'b110, 3'b111, 3'b001, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101,
		3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b001,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b111,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b011, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b011, 3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b110, 3'b101, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b110, 3'b000, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001,
		3'b101, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b000, 3'b111, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b011,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b111, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010,
		3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b101, 3'b001, 3'b010, 3'b010, 3'b000, 3'b010, 3'b000, 3'b001, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b101,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b101, 3'b101, 3'b111, 3'b001, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b011, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b101, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b010, 3'b011, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b101, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b000, 3'b110, 3'b001, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b000, 3'b001, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b111, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011,
		3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b011, 3'b010, 3'b000, 3'b001, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111,
		3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b001, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011,
		3'b001, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110,
		3'b110, 3'b011, 3'b111, 3'b100, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b111, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b011, 3'b001, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b101, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b111, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b011, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b000, 3'b110, 3'b010, 3'b000, 3'b010, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b101, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b111, 3'b000, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b000, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b101, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b110, 3'b010,
		3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b011, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b010, 3'b111, 3'b010, 3'b101, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b001, 3'b111, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b111, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b111, 3'b111, 3'b100,
		3'b011, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b011, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b011, 3'b000, 3'b110, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b101, 3'b110, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b000, 3'b110, 3'b000, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b011, 3'b100, 3'b111, 3'b011,
		3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b011, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011,
		3'b101, 3'b011, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b000,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b001, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b011, 3'b110, 3'b010,
		3'b001, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b001, 3'b110, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b011,
		3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b011, 3'b111, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b101, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b110, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b010, 3'b011, 3'b100, 3'b001,
		3'b001, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b000,
		3'b110, 3'b001, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b001, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b011, 3'b111, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b011, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b111,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b000, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b111, 3'b110, 3'b110, 3'b000, 3'b010, 3'b110, 3'b010, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b011, 3'b111, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b001, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b101, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b111, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b010, 3'b011, 3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b111, 3'b111, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b011, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b011, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b101, 3'b101, 3'b011, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b000, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b010, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b101, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100,
		3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b001, 3'b101, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b111, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b101, 3'b010, 3'b001, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b001, 3'b111, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110,
		3'b011, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b110, 3'b010, 3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b101, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b000, 3'b111, 3'b011, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001,
		3'b011, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b001, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b111, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b011, 3'b101, 3'b010,
		3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b001, 3'b011, 3'b010, 3'b110, 3'b100, 3'b011, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b001, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b001, 3'b011, 3'b010, 3'b001, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b001, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b101, 3'b010, 3'b001, 3'b101, 3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b010, 3'b011, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b011, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000,
		3'b001, 3'b001, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b011, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b101,
		3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b011, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b000,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b101, 3'b101, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b001,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b111, 3'b101, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b101, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110,
		3'b101, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b011, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b111, 3'b010, 3'b000, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b111, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b101, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b110, 3'b111, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b110, 3'b101,
		3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b001, 3'b001, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101,
		3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101, 3'b111, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b001, 3'b101, 3'b001, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b000, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011,
		3'b010, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b000, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b110, 3'b001, 3'b100, 3'b110, 3'b001, 3'b001, 3'b110, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110,
		3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b001, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b101,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b011, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b111, 3'b110, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b101, 3'b000, 3'b110, 3'b001, 3'b000, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b101, 3'b011, 3'b010, 3'b001, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b111, 3'b011, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b101, 3'b111, 3'b110, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b011,
		3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b101, 3'b111, 3'b100, 3'b111, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b011, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b010, 3'b000, 3'b011, 3'b110, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b111, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b000, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b110, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b001, 3'b101, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b000, 3'b101, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b011, 3'b110, 3'b110, 3'b010, 3'b110, 3'b000, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b111, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b101, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b011, 3'b000, 3'b000, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b111, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001,
		3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b001, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b111, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b011, 3'b010, 3'b111,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b111, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b000, 3'b000, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b110, 3'b111,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b101, 3'b010, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b110, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b000, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b110, 3'b011, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b000, 3'b011, 3'b001, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b011,
		3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b101, 3'b100, 3'b110, 3'b110, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001,
		3'b000, 3'b110, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b001, 3'b111, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b101, 3'b001, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110, 3'b101, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b000, 3'b011, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b101, 3'b010, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b110, 3'b110, 3'b010, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b101, 3'b010, 3'b101, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b110, 3'b110, 3'b101, 3'b001, 3'b100, 3'b010, 3'b000, 3'b110, 3'b111, 3'b010, 3'b111, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b110, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b101, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b001, 3'b011, 3'b101, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110, 3'b000, 3'b110, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b101, 3'b001, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b101, 3'b110, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b001, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b101, 3'b001, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b101, 3'b000, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b111, 3'b111, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b001, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b001, 3'b101, 3'b010, 3'b101, 3'b010, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b101, 3'b010,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b011, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b110, 3'b011, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b001, 3'b101, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b001, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b110,
		3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b111, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b010, 3'b111, 3'b111, 3'b110, 3'b001,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b110, 3'b101, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b011,
		3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b101, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b011, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b110, 3'b011, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b101, 3'b010, 3'b101, 3'b000, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b001, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b101, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b000, 3'b011, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b011,
		3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b011, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b001, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b101, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b110, 3'b110, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b111, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b111, 3'b001, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b011, 3'b000, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b000, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010, 3'b011, 3'b010,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110, 3'b101, 3'b001, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b111, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b111, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b101, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b111, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b101, 3'b111, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b101, 3'b111, 3'b000, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b111, 3'b110, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b101,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001, 3'b011, 3'b110, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b000, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b011, 3'b000, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b001, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b011, 3'b011, 3'b001, 3'b010, 3'b101, 3'b010, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b000, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b001, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b101, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b000, 3'b101, 3'b110, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b000, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b010, 3'b101, 3'b101, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b101, 3'b111, 3'b010, 3'b000, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b111, 3'b101, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b011, 3'b110, 3'b101, 3'b101,
		3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b101, 3'b010, 3'b101, 3'b100,
		3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b001, 3'b000, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b000, 3'b111, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b011, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b010, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b110, 3'b111, 3'b110, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b101,
		3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b110, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b111, 3'b111, 3'b101, 3'b101, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b011, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b011, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000,
		3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b101, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b011, 3'b110, 3'b001, 3'b101, 3'b101, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b001, 3'b010, 3'b011, 3'b010, 3'b101, 3'b001, 3'b011, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b011, 3'b011, 3'b010, 3'b001, 3'b000, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b111, 3'b111, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b011, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b101, 3'b000, 3'b101, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b000, 3'b011, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b111,
		3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b001, 3'b101, 3'b010, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b111, 3'b100, 3'b101, 3'b111, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b101, 3'b101, 3'b111,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b001, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b111, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b101, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b011, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b101, 3'b001, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111,
		3'b010, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b000, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b111, 3'b101, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b110, 3'b111, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110,
		3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b110,
		3'b010, 3'b101, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b101,
		3'b101, 3'b011, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b111,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111,
		3'b010, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b001, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b011, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b001, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b000, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b011,
		3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b000, 3'b010, 3'b101, 3'b100, 3'b011, 3'b111, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b101, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b011, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101,
		3'b111, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b000,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100,
		3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b011,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b110, 3'b000,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b000, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b110, 3'b000, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b111, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b001, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b101, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b111, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b011, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b111, 3'b001,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100, 3'b001,
		3'b101, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b011, 3'b000, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b010, 3'b101, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b001, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b011,
		3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b001, 3'b100, 3'b110, 3'b001, 3'b010, 3'b111, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b111, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b001, 3'b010, 3'b101, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b011, 3'b010, 3'b110, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b111, 3'b110, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b111,
		3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b010, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b111, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b001, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b111, 3'b010, 3'b000, 3'b110, 3'b111, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010,
		3'b111, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b111, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100,
		3'b010, 3'b111, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b111, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b010, 3'b001, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b001, 3'b110, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b011, 3'b110, 3'b000, 3'b011, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b000, 3'b001, 3'b101, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b000, 3'b001, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b011, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b111, 3'b001,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b001, 3'b001, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b000,
		3'b110, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b011, 3'b101, 3'b001, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b001, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b111,
		3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b110, 3'b011,
		3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b110, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b101, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b111, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b111,
		3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b011, 3'b110, 3'b010,
		3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b101,
		3'b011, 3'b000, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b000, 3'b010, 3'b001, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b111,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b111, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b011, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b011, 3'b111, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b011, 3'b000, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b011, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b000, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b011, 3'b001, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b000, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b101, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001,
		3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011,
		3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b111, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b000, 3'b101, 3'b001, 3'b010,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b001, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001,
		3'b000, 3'b000, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b101, 3'b001, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110,
		3'b111, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100,
		3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b001, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b001, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b101,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b011, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b111, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b111, 3'b011,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b001, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b111, 3'b001, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b010, 3'b101, 3'b110, 3'b010, 3'b101, 3'b000, 3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b111, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b101, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b101, 3'b110, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b011, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b000, 3'b011,
		3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010,
		3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b010, 3'b110,
		3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b011, 3'b111, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b001, 3'b100, 3'b011,
		3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b101, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b010, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b000, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b101, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b001,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b000, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b000, 3'b000, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b000, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b111, 3'b010, 3'b101, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b111, 3'b110, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b101, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b101, 3'b011, 3'b011, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b010, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b001, 3'b110, 3'b101, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b111, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b011, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b011,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b111, 3'b101, 3'b100, 3'b000,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b111, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b101, 3'b011, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b001, 3'b000, 3'b110, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b101, 3'b010, 3'b001, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b111, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b011, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b001, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b111, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b001, 3'b110, 3'b010,
		3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b001, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b001, 3'b101,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b011, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b001, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b101,
		3'b011, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b110, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b000, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b001, 3'b101, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b000, 3'b110, 3'b001, 3'b011, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b110, 3'b101, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b000, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b110, 3'b110,
		3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b101, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b110, 3'b111, 3'b110,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b011, 3'b010, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101,
		3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b001, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b111, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b101, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b111,
		3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b001, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111,
		3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b000, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001,
		3'b001, 3'b110, 3'b110, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b110, 3'b010, 3'b011, 3'b000, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b000, 3'b111, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b011, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b000, 3'b111, 3'b110, 3'b010, 3'b111, 3'b101, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b111, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b011, 3'b110, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b011, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b001, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b011, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b010, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b000, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b011, 3'b110, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b001, 3'b111, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b111, 3'b101, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b001, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b011, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b011, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b101, 3'b101,
		3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b010, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b101, 3'b111, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b111, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b001, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111,
		3'b011, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b000, 3'b111, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b001,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b001, 3'b110, 3'b011, 3'b010, 3'b011, 3'b010, 3'b111, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b110, 3'b001, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b011,
		3'b001, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b111,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b101, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b111, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b000, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b111, 3'b101, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b110, 3'b000, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b111, 3'b001, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b011,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b101, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b011, 3'b010, 3'b011, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b101,
		3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b011,
		3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b110, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b000, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b101, 3'b001, 3'b101, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b111, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b110, 3'b000, 3'b110, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b101, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b001,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b011,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001,
		3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b000,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b111, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b010, 3'b101, 3'b000, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010,
		3'b001, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011,
		3'b110, 3'b110, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000, 3'b001, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b011, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b101, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000,
		3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b011, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b110, 3'b101, 3'b101,
		3'b100, 3'b111, 3'b110, 3'b000, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b011, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b111, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b110, 3'b101, 3'b110, 3'b011, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b111, 3'b111, 3'b110, 3'b001, 3'b110, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b011, 3'b000,
		3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110,
		3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b111, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b111, 3'b110, 3'b010, 3'b010, 3'b101, 3'b111, 3'b010,
		3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b000, 3'b011, 3'b011, 3'b110, 3'b100, 3'b011,
		3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000,
		3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b100, 3'b000, 3'b111, 3'b000, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b010, 3'b101, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b000, 3'b111, 3'b001, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b001, 3'b011, 3'b110, 3'b011, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b111, 3'b101, 3'b001, 3'b110, 3'b011, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b111, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b000,
		3'b001, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110,
		3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b010, 3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b011, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b011, 3'b001, 3'b010, 3'b111,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b101, 3'b101, 3'b101, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b011, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b000, 3'b001, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b011,
		3'b111, 3'b000, 3'b111, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b101, 3'b110, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111, 3'b001, 3'b000, 3'b010, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b001, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b111, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b011, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b101, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b000, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b011, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b111, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b001, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b001, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b011, 3'b001, 3'b010, 3'b110, 3'b001, 3'b001, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b000, 3'b110, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b111, 3'b101, 3'b100, 3'b010, 3'b110, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b101, 3'b011,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b001, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b001, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b101, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b010, 3'b001, 3'b100, 3'b110, 3'b011, 3'b011, 3'b101, 3'b010, 3'b010, 3'b010, 3'b000, 3'b111, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b001, 3'b011, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110,
		3'b110, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b010, 3'b110, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110,
		3'b110, 3'b011, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b110,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b000, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010,
		3'b111, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b111, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b010, 3'b111, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b010, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b101, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b011, 3'b110, 3'b010, 3'b101, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b000, 3'b010, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b010, 3'b001, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b110, 3'b000,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110,
		3'b111, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010,
		3'b101, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b001, 3'b011, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b001, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b011, 3'b110, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b011, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b010, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b111, 3'b110, 3'b110, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b110, 3'b101, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b010, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b000, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b000, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b001, 3'b100, 3'b101, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b011, 3'b000, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b111, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b011, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b110, 3'b101, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b000, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b011, 3'b001,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b111, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b000, 3'b111, 3'b010, 3'b101, 3'b110, 3'b011, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b110,
		3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b101, 3'b110, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b001, 3'b001, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b101,
		3'b000, 3'b100, 3'b011, 3'b000, 3'b001, 3'b010, 3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b111, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b111, 3'b011, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011,
		3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b101, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b101, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b000, 3'b000, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b011,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b101, 3'b000, 3'b001, 3'b010, 3'b111,
		3'b000, 3'b010, 3'b100, 3'b011, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b000, 3'b011, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b110, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b011, 3'b010, 3'b010, 3'b001, 3'b010, 3'b000, 3'b000, 3'b100, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b011, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b101,
		3'b000, 3'b110, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b000, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b111,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b001, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b010, 3'b000, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b011, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b110, 3'b111,
		3'b100, 3'b110, 3'b110, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b101, 3'b110, 3'b001, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b000, 3'b111, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b011, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b011, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b001,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b000, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b001, 3'b001, 3'b000, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b000, 3'b110, 3'b100, 3'b011,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b101, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b111,
		3'b010, 3'b101, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b101, 3'b000, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b101, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b001, 3'b010, 3'b010, 3'b000, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b010, 3'b111, 3'b111, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b001, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b010, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b110, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b010, 3'b101,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000,
		3'b001, 3'b001, 3'b101, 3'b010, 3'b110, 3'b011, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b000, 3'b101,
		3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b101, 3'b000, 3'b100, 3'b011, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b110, 3'b101,
		3'b110, 3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b101, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b000, 3'b001, 3'b011, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b001,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b011,
		3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b001, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b101, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b000, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b001, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b101,
		3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b001, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011,
		3'b011, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b111, 3'b011, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b111, 3'b110, 3'b110, 3'b001, 3'b100, 3'b110, 3'b001, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b111, 3'b010, 3'b000, 3'b011,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b111, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b101, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b110, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b011, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b000, 3'b001, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b001,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b000,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b000,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110,
		3'b000, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b011, 3'b000, 3'b000, 3'b010, 3'b001, 3'b111,
		3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b001, 3'b011, 3'b010, 3'b111, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b011, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b111, 3'b011, 3'b100, 3'b100, 3'b111, 3'b001, 3'b111, 3'b000, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b000, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b000, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b111, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b101, 3'b110, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b110, 3'b011, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b000, 3'b101, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b000, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010,
		3'b010, 3'b111, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b110,
		3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b010, 3'b000,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b101, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b000, 3'b011, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b101,
		3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001, 3'b011, 3'b111,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011,
		3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b101, 3'b010, 3'b111, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b011, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b011, 3'b000, 3'b011, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b000, 3'b000, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101, 3'b000, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b001, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b101, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b001, 3'b101, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010,
		3'b100, 3'b011, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b001, 3'b010, 3'b111, 3'b100, 3'b000, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b011, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b110, 3'b011, 3'b010, 3'b011, 3'b101,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b111, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b111, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b101, 3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b011, 3'b000, 3'b001, 3'b010,
		3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b001, 3'b111, 3'b111, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b011, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b101, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b001, 3'b101, 3'b100, 3'b000, 3'b010, 3'b000, 3'b011, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b011, 3'b111, 3'b010, 3'b101, 3'b110, 3'b110, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b011, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000,
		3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b001, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b111, 3'b000, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b001, 3'b101, 3'b011, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b101, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b011, 3'b110, 3'b001, 3'b101, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b011, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b010, 3'b001, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b101, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101,
		3'b110, 3'b111, 3'b100, 3'b000, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010,
		3'b101, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b011, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b111, 3'b011, 3'b111, 3'b100, 3'b001, 3'b110, 3'b011, 3'b010, 3'b110, 3'b111, 3'b100, 3'b000,
		3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b101, 3'b001, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b001, 3'b101, 3'b000, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b000, 3'b011, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b011, 3'b100, 3'b010, 3'b111, 3'b111, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b011, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b111, 3'b010, 3'b110,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b011, 3'b000, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b011, 3'b001, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b111, 3'b111, 3'b111, 3'b011, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b011, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b000, 3'b110, 3'b001, 3'b101, 3'b010, 3'b001, 3'b001,
		3'b110, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b111, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b101, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b011, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b000, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b000, 3'b000, 3'b010, 3'b101, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b011, 3'b001, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110,
		3'b001, 3'b001, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b010,
		3'b011, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b011, 3'b110, 3'b010, 3'b000, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b101, 3'b111, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b010, 3'b110,
		3'b110, 3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b111, 3'b111, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b011, 3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b001, 3'b110, 3'b110, 3'b101, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b011,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100,
		3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b011, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b101, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b011, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b000, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b001, 3'b100, 3'b110, 3'b110, 3'b001, 3'b111, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b111, 3'b101, 3'b001,
		3'b010, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b111, 3'b001, 3'b001, 3'b111, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b111, 3'b010, 3'b010,
		3'b111, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b011, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b110, 3'b011, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b011,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101, 3'b111, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b001, 3'b000, 3'b010,
		3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b001, 3'b000, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b000, 3'b010, 3'b111, 3'b101, 3'b010, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b000, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b001, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b101, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b111, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011,
		3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b000, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b010, 3'b001, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b011, 3'b101, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b001, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b110,
		3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b001, 3'b010, 3'b110,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b101, 3'b110, 3'b110, 3'b101, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b001,
		3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b111, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100,
		3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b111, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b101, 3'b101, 3'b101,
		3'b010, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b011, 3'b001, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b111,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b011, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b000, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b111,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b001,
		3'b000, 3'b001, 3'b101, 3'b110, 3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b111, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b111, 3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b111, 3'b001, 3'b101, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b011, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b001, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b101, 3'b100, 3'b001, 3'b001, 3'b101, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b000,
		3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001,
		3'b110, 3'b101, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b001, 3'b110, 3'b000, 3'b101, 3'b100, 3'b111, 3'b101, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b111,
		3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b011, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b111, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b001, 3'b110, 3'b100, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b001, 3'b011, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b101, 3'b011, 3'b110, 3'b001, 3'b110, 3'b010, 3'b011, 3'b010,
		3'b010, 3'b011, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b001, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b111,
		3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b011, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b011, 3'b000, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b111, 3'b110, 3'b100, 3'b000, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b101, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b000, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b001, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001,
		3'b110, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b111, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b111, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b101, 3'b100, 3'b011, 3'b010, 3'b011, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b001,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b110, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b011, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b011, 3'b111, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b000, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b011, 3'b110, 3'b011, 3'b100, 3'b110, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b100, 3'b111, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b110, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b111, 3'b101, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b011, 3'b011, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b000,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b001, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b001, 3'b100, 3'b111, 3'b000, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b010, 3'b111,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b101, 3'b000, 3'b010, 3'b110, 3'b011, 3'b000, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b000, 3'b001, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b010, 3'b011, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b010, 3'b111,
		3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b011, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010,
		3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b111, 3'b001, 3'b100, 3'b010, 3'b110, 3'b101, 3'b111, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b011, 3'b001, 3'b000, 3'b111, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b011, 3'b000, 3'b010, 3'b010, 3'b110, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b010, 3'b000, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b101, 3'b011,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b111, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b010, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b000,
		3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b011, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b011, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b101, 3'b000, 3'b001,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b010, 3'b011, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b000, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b000, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b101, 3'b110, 3'b110, 3'b010, 3'b110, 3'b101, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b011, 3'b000, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110,
		3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110,
		3'b000, 3'b110, 3'b001, 3'b011, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b001, 3'b001, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b000, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b000,
		3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b000, 3'b110, 3'b111, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b001, 3'b101, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b001, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b001, 3'b111, 3'b011, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101,
		3'b011, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b101, 3'b111, 3'b100, 3'b100, 3'b101, 3'b000,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b101, 3'b101, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b101, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b110,
		3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111, 3'b101,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b110, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b000, 3'b001, 3'b101, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b000, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b110, 3'b111, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b110, 3'b000, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b111,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b110, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b000, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b110,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b110, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b110, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111,
		3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b010, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b101, 3'b011, 3'b111, 3'b101, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b011, 3'b000, 3'b000, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b101, 3'b001, 3'b001, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b011, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b010, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b000,
		3'b101, 3'b011, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110, 3'b011, 3'b010, 3'b011, 3'b010, 3'b111, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b000, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b101, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b101,
		3'b111, 3'b010, 3'b111, 3'b101, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b101, 3'b110, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b100, 3'b000, 3'b110, 3'b111, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b000, 3'b001, 3'b000, 3'b101, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b101, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b101, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b110, 3'b010, 3'b111, 3'b001, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b101, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b011, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b011, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b011,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b011, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b000, 3'b101, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100,
		3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b011, 3'b010, 3'b110, 3'b110, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b011, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b001, 3'b011, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b111, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b001, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111,
		3'b110, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b101, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b111, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b111, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b111, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b110, 3'b011, 3'b001, 3'b001, 3'b100, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b000, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b110, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b011,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b011, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b110, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110,
		3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b001, 3'b010, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b111, 3'b111, 3'b010, 3'b000, 3'b010, 3'b001, 3'b010, 3'b001, 3'b001, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b001, 3'b000, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b100, 3'b011, 3'b101, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b001, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b101, 3'b111, 3'b110, 3'b010, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b001,
		3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b111, 3'b111, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b011, 3'b010, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b001, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b000, 3'b000, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b101, 3'b101, 3'b110, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b011, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b001, 3'b101, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b101, 3'b010, 3'b100, 3'b111, 3'b111, 3'b011, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b000, 3'b011, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b111, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b101, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b110, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b010, 3'b111, 3'b010, 3'b101, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b000, 3'b000, 3'b000, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b111, 3'b111, 3'b010, 3'b000, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b111,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b001, 3'b101, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b001, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101,
		3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b011, 3'b111, 3'b010, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b111, 3'b111, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b111,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101,
		3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b000, 3'b010, 3'b101,
		3'b111, 3'b110, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b011, 3'b001, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b011, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b011, 3'b010,
		3'b001, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b101, 3'b010, 3'b111, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b101, 3'b101, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000, 3'b010, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110,
		3'b111, 3'b010, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b111, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b110, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b101, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b011, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b111, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b111, 3'b001, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b111, 3'b001, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b111, 3'b000, 3'b111, 3'b010, 3'b010, 3'b000, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001,
		3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b110, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b001, 3'b001, 3'b111, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b101, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b000, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b000, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b001, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b101,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000,
		3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b011, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b000, 3'b000, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b111, 3'b001,
		3'b001, 3'b010, 3'b000, 3'b110, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b011, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b111, 3'b000, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b011, 3'b111, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b001,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b011, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b011, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111,
		3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b101, 3'b000, 3'b000,
		3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b101, 3'b000, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b010, 3'b011, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b011, 3'b000,
		3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b000, 3'b011, 3'b100, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b010, 3'b101, 3'b001, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b101,
		3'b000, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b110,
		3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b011, 3'b010, 3'b111, 3'b000, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b111, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b111, 3'b001, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b001, 3'b110, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b011, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b101, 3'b110, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b000, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b011, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b000, 3'b110, 3'b101, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010,
		3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b111,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b110, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b101, 3'b000, 3'b100, 3'b110,
		3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b111, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b011, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b110, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b011,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b101, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b110,
		3'b111, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b110, 3'b101, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b011,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b011, 3'b010, 3'b011, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111,
		3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b011, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b000, 3'b110, 3'b011, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b101,
		3'b101, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b000, 3'b000, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b101, 3'b001, 3'b000, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b001, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b001, 3'b000, 3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b111, 3'b011, 3'b000,
		3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b110, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b111, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b011, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b110, 3'b101, 3'b011, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b001, 3'b100, 3'b001, 3'b010, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b101, 3'b101, 3'b100,
		3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b001, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b101, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b010, 3'b010, 3'b001, 3'b000, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010,
		3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b111, 3'b001, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b101, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b111, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b011, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b101, 3'b001, 3'b000, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b101, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b101, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b000, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b110, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b101, 3'b011,
		3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b000,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b111, 3'b100, 3'b010,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b101, 3'b111, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b001,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b111,
		3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b101, 3'b011, 3'b010, 3'b110, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110,
		3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b101, 3'b100, 3'b101, 3'b111, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b001,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b101, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b101, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b101, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b101, 3'b110, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b011, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b011, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b011, 3'b100, 3'b001, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100,
		3'b100, 3'b000, 3'b011, 3'b101, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b111, 3'b000, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b111, 3'b010, 3'b010, 3'b110, 3'b101, 3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b101, 3'b011, 3'b110, 3'b111, 3'b011, 3'b101, 3'b110, 3'b110, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b011, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b000, 3'b010, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b110, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b000, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b011, 3'b011, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b101, 3'b101, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b001, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b000, 3'b101,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b011, 3'b010, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b011, 3'b010, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b001, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b011, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b011, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010,
		3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b111, 3'b011, 3'b111,
		3'b111, 3'b100, 3'b101, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b011, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b110, 3'b010, 3'b011, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b001, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b000, 3'b011,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b110, 3'b001, 3'b001, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b110, 3'b010, 3'b111,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b001, 3'b001, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b010, 3'b011, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b010, 3'b010, 3'b111, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b011, 3'b011, 3'b000,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b000, 3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b000, 3'b100, 3'b111, 3'b101, 3'b101, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b011, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b000, 3'b101, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b000, 3'b011, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b001, 3'b110, 3'b110, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b111, 3'b011, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b000, 3'b111,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b010, 3'b000, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b001,
		3'b011, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b000,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b011, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b101, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b101, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b001, 3'b110, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b110, 3'b001, 3'b000, 3'b100, 3'b101, 3'b010, 3'b111, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b101, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b011, 3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b011, 3'b000, 3'b000, 3'b000, 3'b010, 3'b110,
		3'b000, 3'b001, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110,
		3'b010, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b011, 3'b111, 3'b100, 3'b001, 3'b010, 3'b001,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b110, 3'b010, 3'b011, 3'b111, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b111, 3'b101, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b101, 3'b111, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b101, 3'b010, 3'b111, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b111, 3'b111, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b101, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b101, 3'b010, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b001, 3'b110, 3'b011, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b011, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b111, 3'b000, 3'b010, 3'b001, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b110, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b011, 3'b110, 3'b100, 3'b010, 3'b011, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b001, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b001, 3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b111, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b111,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b000, 3'b100, 3'b111, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b011, 3'b000, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b000, 3'b010, 3'b000,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b111, 3'b110, 3'b011, 3'b001, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b110, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b111, 3'b101, 3'b011, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b011, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b110, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b011, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b111, 3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b101, 3'b101, 3'b111, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b101,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b001, 3'b100, 3'b000, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b110, 3'b110, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b000, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b101, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b011, 3'b111,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b111, 3'b010, 3'b111, 3'b000, 3'b100, 3'b011, 3'b000, 3'b010, 3'b010, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b001, 3'b110, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b000, 3'b100, 3'b010, 3'b011, 3'b010, 3'b101, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b000, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011,
		3'b001, 3'b000, 3'b010, 3'b000, 3'b010, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b110, 3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b101, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b101, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b011, 3'b011, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b101, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b001, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b001, 3'b001, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b110, 3'b011, 3'b110, 3'b010,
		3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b110, 3'b000, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b011, 3'b111, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b101,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b111,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b101, 3'b110, 3'b101, 3'b100, 3'b001,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b101, 3'b001, 3'b000, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b010, 3'b000, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b000, 3'b110, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b001, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b010, 3'b101, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b010,
		3'b000, 3'b011, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b001,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101,
		3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b110, 3'b010, 3'b001, 3'b011, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b101, 3'b001, 3'b010, 3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b110, 3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b101, 3'b011, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b101, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b111, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b111, 3'b000, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b110,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b101, 3'b111, 3'b010, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b101, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010,
		3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b001, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b010, 3'b000, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b011, 3'b000, 3'b001,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b011, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b110, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b111, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b011, 3'b010, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b101,
		3'b001, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b000, 3'b000, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110, 3'b010, 3'b000, 3'b011, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b000, 3'b101, 3'b100, 3'b101, 3'b010, 3'b001, 3'b011, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b011, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b011, 3'b010, 3'b101, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b111,
		3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b101, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111, 3'b000, 3'b000, 3'b100, 3'b001, 3'b010, 3'b001,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b101, 3'b000, 3'b001, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b001, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b010, 3'b101, 3'b010, 3'b111,
		3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b000, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b011, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b111, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b000,
		3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b001, 3'b111, 3'b110, 3'b101, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b110, 3'b000, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b000, 3'b100, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b001, 3'b001, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110,
		3'b111, 3'b000, 3'b111, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b010, 3'b001, 3'b111, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b000, 3'b101, 3'b001,
		3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b001, 3'b011, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b000, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b001, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b000, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b010, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b000, 3'b010, 3'b000, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b111, 3'b111, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b110,
		3'b011, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b101, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b101, 3'b010, 3'b000, 3'b000, 3'b011, 3'b010, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010,
		3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b011, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b001,
		3'b001, 3'b100, 3'b010, 3'b011, 3'b001, 3'b011, 3'b110, 3'b010, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b110, 3'b001, 3'b000, 3'b100, 3'b110, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b001,
		3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b011, 3'b011, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b101, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b101, 3'b000, 3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b000, 3'b100, 3'b011,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b000, 3'b001, 3'b111, 3'b001, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b101, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b001, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b011, 3'b111, 3'b100, 3'b010,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b011, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b110, 3'b100, 3'b111, 3'b010, 3'b011, 3'b000,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b000, 3'b010, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000,
		3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b111, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b111, 3'b100, 3'b011, 3'b001,
		3'b010, 3'b000, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b111, 3'b110, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b111, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111, 3'b110, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b111, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b111, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b011, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b000, 3'b101, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b011,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b011, 3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b101, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b111, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b110, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b011, 3'b100, 3'b101, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b101, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b000, 3'b100, 3'b010, 3'b000, 3'b001, 3'b010, 3'b001, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110,
		3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b111, 3'b100, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b110, 3'b111, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b111, 3'b101, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000,
		3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b110, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b011, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b001, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110,
		3'b101, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110,
		3'b010, 3'b011, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b111, 3'b010, 3'b011, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b001, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b011, 3'b101, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b011, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b101, 3'b011, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b010, 3'b000, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b110, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b001, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b001, 3'b101, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b111, 3'b110,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110,
		3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b110, 3'b111, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b000, 3'b101, 3'b011, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b101, 3'b101, 3'b010,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010,
		3'b110, 3'b000, 3'b101, 3'b000, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b000, 3'b001, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b001, 3'b111,
		3'b011, 3'b010, 3'b000, 3'b000, 3'b101, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000, 3'b101, 3'b101, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b111, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b001, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b010, 3'b101, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b000, 3'b111, 3'b011, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b011, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b011, 3'b000, 3'b100, 3'b011, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b101, 3'b110, 3'b001, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b110, 3'b010, 3'b110, 3'b110, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b011, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b111, 3'b011,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b110, 3'b010, 3'b110, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b111, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b011, 3'b100, 3'b000, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b111, 3'b100, 3'b000, 3'b010,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b101, 3'b001, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b001, 3'b010, 3'b111, 3'b111, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b011, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b011, 3'b101, 3'b100, 3'b001, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b010, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b000, 3'b101, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b011, 3'b101, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b110, 3'b011, 3'b100, 3'b101, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101,
		3'b110, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b011,
		3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b111, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b001, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b110,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000, 3'b011, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b101, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b011,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b111, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b000, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b110, 3'b001, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b000, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b011, 3'b110, 3'b011, 3'b100, 3'b000, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b011, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b101, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b101,
		3'b100, 3'b100, 3'b000, 3'b111, 3'b111, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b110, 3'b001, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b101, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b111, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b111, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101,
		3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b111, 3'b000, 3'b001, 3'b101, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b111, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b101, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b111, 3'b100, 3'b110, 3'b101, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b101, 3'b111, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b011,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110, 3'b001, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b101,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b111, 3'b101, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000,
		3'b000, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b011, 3'b001,
		3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b110, 3'b101, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b010, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b011,
		3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110,
		3'b011, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b000, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001, 3'b110, 3'b100,
		3'b001, 3'b000, 3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b111, 3'b001, 3'b000, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b001, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b101, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b011, 3'b101, 3'b011, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b011, 3'b010, 3'b100, 3'b000, 3'b011,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b010, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b101, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b011, 3'b101, 3'b010, 3'b000, 3'b011, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b001, 3'b110, 3'b001, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b101, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b101, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b101, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b001, 3'b100, 3'b110, 3'b001, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b110, 3'b111, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b010, 3'b111, 3'b101, 3'b110, 3'b110, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b101, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b000, 3'b000,
		3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b111, 3'b010,
		3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b111, 3'b011, 3'b110, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b000, 3'b010, 3'b001, 3'b110, 3'b100, 3'b001,
		3'b011, 3'b001, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000,
		3'b100, 3'b101, 3'b010, 3'b000, 3'b001, 3'b101, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b111, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b011, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b000, 3'b111, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000,
		3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b010, 3'b111, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b001,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b111, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b111,
		3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b101, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b011, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100,
		3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b011, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b001, 3'b111, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b010, 3'b000, 3'b001,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b011, 3'b010, 3'b011, 3'b100, 3'b000, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b111,
		3'b110, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b000, 3'b001, 3'b101, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000,
		3'b010, 3'b000, 3'b011, 3'b000, 3'b010, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b111, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b011, 3'b000, 3'b100, 3'b011, 3'b010, 3'b101, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b000, 3'b011, 3'b011, 3'b111, 3'b101, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b011, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b011, 3'b110, 3'b010, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b101, 3'b001, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b101, 3'b000, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b101, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b111, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b011, 3'b101,
		3'b101, 3'b101, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b011, 3'b100, 3'b110, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000,
		3'b001, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b000, 3'b001, 3'b010, 3'b000, 3'b001, 3'b111, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b101,
		3'b111, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b111,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b011, 3'b000, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b101, 3'b001, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b011, 3'b110, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b101, 3'b011, 3'b010, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b011, 3'b010, 3'b011,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b011, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b111,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b111, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111,
		3'b101, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b111, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b100, 3'b011, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b111, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b101,
		3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b110,
		3'b110, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100,
		3'b110, 3'b111, 3'b110, 3'b110, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b011, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b111, 3'b100,
		3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b101, 3'b010, 3'b110, 3'b111, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b000, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b011, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b001, 3'b011, 3'b101,
		3'b010, 3'b100, 3'b111, 3'b001, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b110, 3'b000, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b000, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b011, 3'b100, 3'b101, 3'b000, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b111, 3'b101, 3'b000, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b111,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b000, 3'b011, 3'b000, 3'b100, 3'b101, 3'b010, 3'b110, 3'b000, 3'b001, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b010, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b111,
		3'b100, 3'b011, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001, 3'b010, 3'b001, 3'b110, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b111,
		3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b111, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b010,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b011, 3'b001, 3'b100, 3'b011, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b101, 3'b100, 3'b111, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b000, 3'b111, 3'b001, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b000, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b000, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b101, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b111, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b010, 3'b101, 3'b011, 3'b100, 3'b111, 3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b000, 3'b111, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b000, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b101, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b110, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b001, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b011, 3'b001, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b101, 3'b100, 3'b000, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101,
		3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b110, 3'b010,
		3'b000, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b000, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b010, 3'b010, 3'b010, 3'b111, 3'b111, 3'b100, 3'b010, 3'b111, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b111, 3'b110, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b011, 3'b001, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b011, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b011, 3'b000, 3'b111, 3'b111, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100,
		3'b011, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b101, 3'b001, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b111, 3'b110, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b011, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001,
		3'b001, 3'b101, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b111, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b001, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100, 3'b001, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b100, 3'b111, 3'b110, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110, 3'b101, 3'b101, 3'b100, 3'b100, 3'b101, 3'b010, 3'b001, 3'b100, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b111, 3'b110,
		3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b011, 3'b011, 3'b101, 3'b001, 3'b110,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b101, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b000, 3'b000, 3'b100,
		3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b110, 3'b010, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b100, 3'b110, 3'b100, 3'b000, 3'b111, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101,
		3'b110, 3'b110, 3'b101, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b010,
		3'b101, 3'b111, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b101, 3'b010, 3'b111, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b000, 3'b010, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b101, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b110, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b000, 3'b011, 3'b110, 3'b001,
		3'b100, 3'b110, 3'b100, 3'b101, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b001, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b000, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b000, 3'b001, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001,
		3'b110, 3'b101, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010, 3'b011, 3'b101, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b011, 3'b110, 3'b100, 3'b010, 3'b101, 3'b010, 3'b001, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b100, 3'b011, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b000, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b101, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b001, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b000, 3'b110, 3'b111, 3'b010, 3'b111, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b110, 3'b000, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b001, 3'b011, 3'b001, 3'b111, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b000, 3'b001, 3'b010, 3'b110, 3'b011,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b011, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b101, 3'b010, 3'b111, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b000, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000, 3'b011,
		3'b010, 3'b011, 3'b010, 3'b011, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b001, 3'b110, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b000, 3'b111, 3'b011, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b000,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b001, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b110, 3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b000, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b110, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b110, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111,
		3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b110, 3'b100, 3'b011, 3'b111, 3'b110, 3'b001, 3'b100,
		3'b000, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b110, 3'b100, 3'b110, 3'b110, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b111, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b110, 3'b110, 3'b110, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b001, 3'b100, 3'b110, 3'b011, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b001,
		3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b000, 3'b100, 3'b010, 3'b110, 3'b111, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b111, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b001,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b110, 3'b010, 3'b010, 3'b110, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b011, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b111, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101,
		3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b011, 3'b110,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b111, 3'b101, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b011, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b010, 3'b001, 3'b010, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011,
		3'b101, 3'b001, 3'b000, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b010, 3'b011, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b111, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b111, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b000, 3'b111, 3'b000, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b101, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b101, 3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b000, 3'b010, 3'b011,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b101, 3'b100, 3'b111, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b010, 3'b110, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b000, 3'b100, 3'b010, 3'b110, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b000, 3'b100, 3'b000, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010,
		3'b011, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b111, 3'b000, 3'b100, 3'b110, 3'b100, 3'b101, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b010, 3'b010, 3'b111, 3'b001, 3'b010, 3'b000, 3'b000,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b000, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b101, 3'b011, 3'b000, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b001, 3'b101, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b001, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b010, 3'b001, 3'b010, 3'b110, 3'b011, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b000, 3'b010, 3'b100,
		3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b000, 3'b101, 3'b101, 3'b100, 3'b110, 3'b110, 3'b001,
		3'b111, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b110, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b000, 3'b110, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b000, 3'b101,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b000, 3'b000,
		3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110,
		3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b110,
		3'b010, 3'b100, 3'b000, 3'b010, 3'b011, 3'b111, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b000, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b000, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100,
		3'b010, 3'b101, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b011, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b011, 3'b011, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b111, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b101, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b101, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b110, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b111, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b111, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b110, 3'b010, 3'b000, 3'b101, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b000, 3'b110, 3'b111, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b010, 3'b100, 3'b010, 3'b011, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b000, 3'b101, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b011, 3'b000, 3'b100, 3'b110, 3'b111, 3'b010, 3'b110, 3'b010,
		3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b011, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b111, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b000, 3'b001, 3'b001, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b010, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b001, 3'b011, 3'b111, 3'b110, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110,
		3'b000, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b101, 3'b010, 3'b100, 3'b000, 3'b111, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b111, 3'b001, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b000, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b111,
		3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b101, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b001, 3'b110, 3'b101, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b111, 3'b011, 3'b101, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b001, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b101, 3'b100, 3'b011, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b000, 3'b010, 3'b101, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b011, 3'b100, 3'b001, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b101, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b000, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b000, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b000, 3'b100, 3'b011, 3'b000, 3'b101, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111,
		3'b110, 3'b110, 3'b100, 3'b001, 3'b011, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b010, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b001, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b111, 3'b000, 3'b101, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b000, 3'b010, 3'b100, 3'b011, 3'b110, 3'b100, 3'b101, 3'b000, 3'b011, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b101, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b110, 3'b011, 3'b101, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b011, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b101, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b000, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b000, 3'b101, 3'b110, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b101, 3'b010, 3'b000, 3'b100, 3'b110, 3'b001, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b011, 3'b101, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b111, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b010, 3'b011, 3'b100, 3'b100, 3'b111, 3'b000, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b111, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b010,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100,
		3'b010, 3'b111, 3'b111, 3'b011, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b011, 3'b010, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b111, 3'b111, 3'b100, 3'b100, 3'b000, 3'b101, 3'b010, 3'b010, 3'b001, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b000, 3'b110, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b000, 3'b100, 3'b011,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b000, 3'b000, 3'b101, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111, 3'b101, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b011, 3'b001,
		3'b110, 3'b100, 3'b111, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b110, 3'b100, 3'b001, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b110, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b001,
		3'b101, 3'b100, 3'b000, 3'b101, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b101, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b110, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b001, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b101, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b011, 3'b110, 3'b010, 3'b100, 3'b001, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b010, 3'b000,
		3'b011, 3'b011, 3'b100, 3'b010, 3'b001, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b011, 3'b100, 3'b101, 3'b100, 3'b111, 3'b001, 3'b110, 3'b010, 3'b000, 3'b111,
		3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b010, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b111, 3'b111, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b101, 3'b000, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b011, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b110, 3'b000, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010,
		3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b000,
		3'b100, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b001, 3'b111, 3'b100, 3'b001, 3'b010, 3'b001, 3'b001, 3'b110, 3'b010, 3'b101, 3'b110, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b011, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b100, 3'b110, 3'b011, 3'b110, 3'b110, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b110, 3'b100, 3'b000, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010,
		3'b010, 3'b001, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b011, 3'b001, 3'b010, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b001, 3'b100, 3'b110,
		3'b101, 3'b110, 3'b111, 3'b100, 3'b111, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b001, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110,
		3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b000,
		3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b010, 3'b110, 3'b100, 3'b011, 3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b100, 3'b011, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b001, 3'b010, 3'b101, 3'b111, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b101, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b010, 3'b110, 3'b110, 3'b100, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b000, 3'b111, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b111, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010,
		3'b110, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b100, 3'b100, 3'b000, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b001, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b000, 3'b000, 3'b000, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b110, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b011, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b101, 3'b000, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b011, 3'b110, 3'b110, 3'b001, 3'b110, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b111, 3'b100, 3'b001, 3'b001,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b000, 3'b011,
		3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010,
		3'b110, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b011, 3'b001, 3'b111, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b101, 3'b100, 3'b001, 3'b111, 3'b100, 3'b101,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b001, 3'b110, 3'b001, 3'b111, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b001,
		3'b001, 3'b001, 3'b110, 3'b101, 3'b110, 3'b100, 3'b011, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b101, 3'b010, 3'b010,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b011, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b111, 3'b111, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b011, 3'b010, 3'b010, 3'b010, 3'b011, 3'b100, 3'b110, 3'b100, 3'b000, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110, 3'b011, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b101, 3'b111, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b011, 3'b010, 3'b100, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b111, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b011, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b101, 3'b110, 3'b110, 3'b010, 3'b101, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b101, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b000, 3'b110, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100,
		3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b111, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b101, 3'b010,
		3'b111, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b101, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b111, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b110, 3'b011, 3'b010, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b001, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b100, 3'b111, 3'b010, 3'b111, 3'b101, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b010, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b011,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b100, 3'b001, 3'b000, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b111,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b001, 3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b101, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b011, 3'b110, 3'b001, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b111, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010, 3'b111, 3'b011, 3'b111, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b011, 3'b010, 3'b100, 3'b101, 3'b000,
		3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b011,
		3'b010, 3'b000, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b001, 3'b010, 3'b110, 3'b001,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110,
		3'b011, 3'b101, 3'b110, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b110, 3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b001, 3'b110, 3'b110, 3'b010, 3'b010, 3'b111, 3'b011, 3'b111, 3'b111, 3'b100, 3'b100, 3'b011, 3'b100,
		3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b011, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b111, 3'b110, 3'b100, 3'b000, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b100, 3'b010, 3'b110, 3'b111, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b001, 3'b011, 3'b100, 3'b100, 3'b001, 3'b100, 3'b011, 3'b101, 3'b010, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b010, 3'b011, 3'b010, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b111, 3'b100,
		3'b001, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100,
		3'b000, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b101, 3'b001, 3'b011, 3'b111, 3'b110, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b011, 3'b100,
		3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b011, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010, 3'b001,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b011, 3'b100, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b110, 3'b111, 3'b100, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b110, 3'b011, 3'b010, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b011, 3'b110, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b011, 3'b100, 3'b111, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b001, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b100,
		3'b110, 3'b001, 3'b010, 3'b111, 3'b010, 3'b100, 3'b101, 3'b101, 3'b010, 3'b100, 3'b001, 3'b111, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001,
		3'b110, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b000, 3'b100, 3'b110, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b100, 3'b101, 3'b000, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110,
		3'b011, 3'b010, 3'b110, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b111, 3'b110, 3'b100, 3'b100, 3'b010, 3'b001, 3'b101, 3'b010, 3'b110, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b111, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b111, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b101,
		3'b010, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b100, 3'b010,
		3'b010, 3'b011, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b110, 3'b011, 3'b010, 3'b110, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b010, 3'b101, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100,
		3'b001, 3'b100, 3'b000, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b110, 3'b111, 3'b100, 3'b110, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b011, 3'b100,
		3'b111, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b010, 3'b001, 3'b100,
		3'b011, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100,
		3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b010, 3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b000,
		3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b001, 3'b100, 3'b010, 3'b111, 3'b001, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b001, 3'b011,
		3'b010, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b110, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b011, 3'b100, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100,
		3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b101, 3'b000, 3'b100, 3'b000, 3'b111,
		3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b110,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b111, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b001, 3'b110, 3'b010, 3'b111, 3'b010, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b110, 3'b010, 3'b011, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b010, 3'b010, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b010, 3'b101, 3'b000, 3'b010, 3'b010, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b011, 3'b001, 3'b010, 3'b000, 3'b010, 3'b010, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b000, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110, 3'b001,
		3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b001, 3'b100, 3'b100, 3'b110, 3'b010,
		3'b111, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b111, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b101, 3'b100, 3'b110, 3'b100, 3'b000, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b001,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b110, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b010, 3'b000, 3'b111, 3'b010, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100,
		3'b001, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b101, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b011, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100,
		3'b111, 3'b100, 3'b001, 3'b100, 3'b101, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b111, 3'b010, 3'b000, 3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b111,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b001, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b110, 3'b000,
		3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b000, 3'b101, 3'b100, 3'b100, 3'b000,
		3'b110, 3'b001, 3'b110, 3'b110, 3'b010, 3'b100, 3'b100, 3'b011, 3'b010, 3'b001, 3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b001, 3'b010, 3'b110, 3'b000, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b001, 3'b100, 3'b111, 3'b110, 3'b110, 3'b100, 3'b111, 3'b110, 3'b011, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b110, 3'b011, 3'b100, 3'b110, 3'b000, 3'b011, 3'b111, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010,
		3'b011, 3'b010, 3'b110, 3'b000, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b101, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b010, 3'b010, 3'b010, 3'b110, 3'b100,
		3'b100, 3'b010, 3'b110, 3'b010, 3'b101, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b001, 3'b110, 3'b110, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b101, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b110, 3'b110, 3'b100, 3'b110, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b101, 3'b010, 3'b110, 3'b000, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b111, 3'b000, 3'b101, 3'b101, 3'b110, 3'b010, 3'b000, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100,
		3'b111, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b010, 3'b110, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100,
		3'b010, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b101, 3'b100,
		3'b000, 3'b111, 3'b001, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b111, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b011, 3'b000, 3'b110, 3'b000, 3'b100,
		3'b011, 3'b101, 3'b110, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b101, 3'b110, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b000, 3'b001, 3'b110, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b011, 3'b111,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100, 3'b101, 3'b100,
		3'b010, 3'b010, 3'b000, 3'b100, 3'b111, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010,
		3'b000, 3'b100, 3'b110, 3'b100, 3'b010, 3'b101, 3'b110, 3'b010, 3'b010, 3'b110, 3'b100, 3'b011, 3'b011, 3'b010, 3'b010, 3'b110, 3'b110, 3'b010, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b111, 3'b100, 3'b110, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b001,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b000, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b001, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100,
		3'b001, 3'b001, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b001, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101,
		3'b110, 3'b001, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b011, 3'b111, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b101, 3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b010, 3'b100, 3'b001, 3'b100, 3'b011, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b110, 3'b100, 3'b111, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b010, 3'b101, 3'b100, 3'b101, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001, 3'b001, 3'b010, 3'b100, 3'b000, 3'b000,
		3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b101, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b101, 3'b010, 3'b100, 3'b110, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b010, 3'b100, 3'b001, 3'b010,
		3'b100, 3'b011, 3'b010, 3'b101, 3'b100, 3'b010, 3'b001, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b110, 3'b010, 3'b101, 3'b100, 3'b010, 3'b011, 3'b100, 3'b010, 3'b111, 3'b010, 3'b100, 3'b110, 3'b010, 3'b001, 3'b110,
		3'b100, 3'b011, 3'b110, 3'b110, 3'b100, 3'b111, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b100, 3'b000, 3'b111, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b000, 3'b110, 3'b001, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b000, 3'b110, 3'b000, 3'b010, 3'b110, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b001, 3'b110, 3'b001, 3'b100, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b111, 3'b100, 3'b010, 3'b001, 3'b110, 3'b111,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b000, 3'b001, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b110, 3'b001, 3'b100, 3'b100, 3'b010, 3'b110, 3'b001, 3'b111, 3'b110, 3'b010, 3'b110, 3'b010, 3'b101,
		3'b100, 3'b001, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b110, 3'b001, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b101, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b001, 3'b101,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b100, 3'b011, 3'b010, 3'b011, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b111, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110,
		3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b110, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b110, 3'b010, 3'b000, 3'b100, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b110, 3'b110, 3'b100,
		3'b110, 3'b000, 3'b010, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b011, 3'b010, 3'b000, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b110, 3'b000, 3'b000, 3'b001, 3'b100, 3'b010, 3'b101, 3'b100, 3'b010, 3'b010,
		3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b010, 3'b001,
		3'b010, 3'b001, 3'b000, 3'b111, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101,
		3'b010, 3'b111, 3'b110, 3'b110, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b010, 3'b010, 3'b110, 3'b101, 3'b100, 3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b101, 3'b010, 3'b100, 3'b100, 3'b001, 3'b001,
		3'b110, 3'b100, 3'b100, 3'b101, 3'b101, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b101, 3'b010, 3'b100, 3'b111, 3'b010, 3'b100, 3'b000, 3'b100, 3'b111, 3'b010, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b001, 3'b000, 3'b100, 3'b100,
		3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b110, 3'b000, 3'b100, 3'b100,
		3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b010, 3'b011, 3'b011, 3'b101, 3'b100, 3'b100, 3'b001, 3'b110, 3'b100, 3'b010, 3'b000, 3'b100, 3'b110,
		3'b000, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b000, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b010, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b100, 3'b110, 3'b000, 3'b101, 3'b111, 3'b110, 3'b100, 3'b101,
		3'b100, 3'b010, 3'b110, 3'b100, 3'b000, 3'b100, 3'b110, 3'b001, 3'b101, 3'b100, 3'b000, 3'b100, 3'b100, 3'b111, 3'b011, 3'b010, 3'b100, 3'b110, 3'b100, 3'b010,
		3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b000, 3'b001, 3'b100, 3'b101, 3'b111, 3'b000, 3'b010, 3'b001, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b110,
		3'b010, 3'b010, 3'b111, 3'b010, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b110, 3'b100, 3'b000, 3'b100, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010,
		3'b100, 3'b100, 3'b110, 3'b000, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b010, 3'b100, 3'b001, 3'b010, 3'b110,
		3'b101, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b010, 3'b100,
		3'b010, 3'b100, 3'b010, 3'b101, 3'b100, 3'b100, 3'b100, 3'b000, 3'b110, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b000, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b011, 3'b100, 3'b011, 3'b010, 3'b010, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b010, 3'b100, 3'b000,
		3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b010, 3'b111, 3'b101, 3'b100, 3'b110, 3'b100, 3'b010, 3'b010, 3'b001, 3'b100, 3'b010, 3'b100, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100,
		3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100, 3'b110, 3'b100, 3'b101, 3'b111, 3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b110, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b010, 3'b011, 3'b100, 3'b011, 3'b000, 3'b100, 3'b001, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b010, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b100, 3'b101, 3'b110, 3'b100, 3'b010, 3'b111, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010,
		3'b001, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b001, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b000, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b001, 3'b110,
		3'b101, 3'b110, 3'b100, 3'b010, 3'b000, 3'b111, 3'b100, 3'b011, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b011, 3'b010, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b110, 3'b100, 3'b100, 3'b100, 3'b001, 3'b100, 3'b001, 3'b110, 3'b000, 3'b010, 3'b100, 3'b110, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b100, 3'b010, 3'b111, 3'b110, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010,
		3'b100, 3'b001, 3'b100, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b110, 3'b110, 3'b110, 3'b011, 3'b100, 3'b110, 3'b100, 3'b100, 3'b001, 3'b010, 3'b100, 3'b110,
		3'b100, 3'b100, 3'b110, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b100, 3'b100, 3'b011, 3'b100, 3'b100, 3'b111, 3'b100, 3'b101, 3'b100, 3'b100,
		3'b100, 3'b010, 3'b100, 3'b110, 3'b100, 3'b011, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b101, 3'b000, 3'b100, 3'b100,
		3'b100, 3'b110, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b010, 3'b100, 3'b110, 3'b110, 3'b101, 3'b010, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100,
		3'b010, 3'b100, 3'b100, 3'b101, 3'b100, 3'b010, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b110, 3'b010,
		3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b101, 3'b110, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b011, 3'b100,
		3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b000, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b000, 3'b010,
		3'b100, 3'b100, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b110, 3'b100, 3'b010, 3'b100, 3'b110,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b111, 3'b010, 3'b010, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b011, 3'b001, 3'b100, 3'b001, 3'b110, 3'b010, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b111, 3'b100, 3'b010, 3'b110, 3'b101, 3'b100, 3'b100, 3'b100, 3'b101, 3'b011, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b101, 3'b100,
		3'b110, 3'b110, 3'b011, 3'b000, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b100, 3'b010, 3'b111, 3'b100, 3'b100, 3'b100, 3'b100, 3'b110, 3'b100,
		3'b001, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 3'b010, 3'b010, 3'b100, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b110,
		3'b111, 3'b110, 3'b100, 3'b110, 3'b001, 3'b110, 3'b100, 3'b100, 3'b100, 3'b100, 3'b101, 3'b001, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100,
		3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b010, 3'b000, 3'b100, 3'b100, 3'b010, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b010,
		3'b101, 3'b110, 3'b001, 3'b010, 3'b100, 3'b011, 3'b001, 3'b110, 3'b100, 3'b100, 3'b000, 3'b011, 3'b100, 3'b110, 3'b111, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100,
		3'b110, 3'b100, 3'b010, 3'b101, 3'b101, 3'b001, 3'b000, 3'b110, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b100, 3'b100, 3'b010, 3'b100, 3'b101, 3'b100, 3'b010
	};
