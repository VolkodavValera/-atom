logic [31:0] Bit_Avalon [12] =
		'{	32'h4334_0000, // 180
			32'h42B4_0000, // 90
			32'h4234_0000, // 45
			32'h41B4_0000, // 22.5
			32'h4134_0000, // 11.25
			32'h40B4_0000, // 5.625
			32'h4034_0000, // 2.8125
			32'h3FB3_F7CE, // 1.4062
			32'h3F33_F7CE, // 0.7031
			32'h3EB3_F7CC, // 0.3516
			32'h3E34_3958, // 0.1758
			32'h3DB4_3950  // 0.0878
		};

logic [31:0] Whole_corners [0:199] =
		'{	32'h0000_0000, 32'h3F66_6666, 32'h3FE6_6666, 32'h402C_CCCC, 32'h4066_6666, 32'h4090_0000, 32'h40AC_CCCC, 32'h40C9_9999, 32'h40E6_6666, 32'h4101_9999,	// 0-8.1
			32'h4110_0000, 32'h411E_6666, 32'h412C_CCCC, 32'h413B_3333, 32'h4149_9999, 32'h4158_0000, 32'h4166_6666, 32'h4174_CCCC, 32'h4181_9999, 32'h4188_CCCC,	// 9-17.1
			32'h4190_0000, 32'h4197_3333, 32'h419E_6666, 32'h41A5_9999, 32'h41AC_CCCC, 32'h41B4_0000, 32'h41BB_3333, 32'h41C2_6666, 32'h41C9_9999, 32'h41D0_CCCC,	// 18-26.1
			32'h41D8_0000, 32'h41DF_3333, 32'h41E6_6666, 32'h41ED_9999, 32'h41F4_CCCC, 32'h41FC_0000, 32'h4201_9999, 32'h4205_3333, 32'h4208_CCCC, 32'h420C_6666,	// 27-35.1
			32'h4210_0000, 32'h4213_9999, 32'h4217_3333, 32'h421A_CCCC, 32'h421E_6666, 32'h4222_0000, 32'h4225_9999, 32'h4229_3333, 32'h422C_CCCC, 32'h4230_6666,	// 36-44.1
			32'h4234_0000, 32'h4237_9999, 32'h423B_3333, 32'h423E_CCCC, 32'h4242_6666, 32'h4246_0000, 32'h4249_9999, 32'h424D_3333, 32'h4250_CCCC, 32'h4254_6666,	// 45-53.1
			32'h4258_0000, 32'h425B_9999, 32'h425F_3333, 32'h4262_CCCC, 32'h4266_6666, 32'h426A_0000, 32'h426D_9999, 32'h4271_3333, 32'h4274_CCCC, 32'h4278_6666,	// 54-62.1
			32'h427C_0000, 32'h427F_9999, 32'h4281_9999, 32'h4283_6666, 32'h4285_3333, 32'h4287_0000, 32'h4288_CCCC, 32'h428A_9999, 32'h428C_6666, 32'h428E_3333,	// 63-71.1
			32'h4290_0000, 32'h4291_CCCC, 32'h4293_9999, 32'h4295_6666, 32'h4297_3333, 32'h4299_0000, 32'h429A_CCCC, 32'h429C_9999, 32'h429E_6666, 32'h42A0_3333,	// 72-80.1
			32'h42A2_0000, 32'h42A3_CCCC, 32'h42A5_9999, 32'h42A7_6666, 32'h42A9_3333, 32'h42AB_0000, 32'h42AC_CCCC, 32'h42AE_9999, 32'h42B0_6666, 32'h42B2_3333, 	// 81-89.1
			32'h42B4_0000, 32'h42B5_CCCC, 32'h42B7_9999, 32'h42B9_6666, 32'h42BB_3333, 32'h42BD_0000, 32'h42BE_CCCC, 32'h42C0_9999, 32'h42C2_6666, 32'h42C4_3333, 	// 90-98.1
			32'h42C6_0000, 32'h42C7_CCCC, 32'h42C9_9999, 32'h42CB_6666, 32'h42CD_3333, 32'h42CF_0000, 32'h42D0_CCCC, 32'h42D2_9999, 32'h42D4_6666, 32'h42D6_3333, 	// 99-107.1
			32'h42D8_0000, 32'h42D9_CCCC, 32'h42DB_9999, 32'h42DD_6666, 32'h42DF_3333, 32'h42E1_0000, 32'h42E2_CCCC, 32'h42E4_9999, 32'h42E6_6666, 32'h42E8_3333, 	// 108-116.1
			32'h42EA_0000, 32'h42EB_CCCC, 32'h42ED_9999, 32'h42EF_6666, 32'h42F1_3333, 32'h42F3_0000, 32'h42F4_CCCC, 32'h42F6_9999, 32'h42F8_6666, 32'h42FA_3333, 	// 117-125.1
			32'h42FC_0000, 32'h42FD_CCCC, 32'h42FF_9999, 32'h4300_B333, 32'h4301_9999, 32'h4302_8000, 32'h4303_6666, 32'h4304_4CCC, 32'h4305_3333, 32'h4306_1999,	// 126-134.1
			32'h4307_0000, 32'h4307_E666, 32'h4308_CCCC, 32'h4309_B333, 32'h430A_9999, 32'h430B_8000, 32'h430C_6666, 32'h430D_4CCC, 32'h430E_3333, 32'h430F_1999, 	// 135-143.1
			32'h4310_0000, 32'h4310_E666, 32'h4311_CCCC, 32'h4312_B333, 32'h4313_9999, 32'h4314_8000, 32'h4315_6666, 32'h4316_4CCC, 32'h4317_3333, 32'h4318_1999, 	// 144-152.1
			32'h4319_0000, 32'h4319_E666, 32'h431A_CCCC, 32'h431B_B333, 32'h431C_9999, 32'h431D_8000, 32'h431E_6666, 32'h431F_4CCC, 32'h4320_3333, 32'h4321_1999,	// 153-161.1
			32'h4322_0000, 32'h4322_E666, 32'h4323_CCCC, 32'h4324_B333, 32'h4325_9999, 32'h4326_8000, 32'h4327_6666, 32'h4328_4CCC, 32'h4329_3333, 32'h432A_1999,	// 162-170.1
			32'h432B_0000, 32'h432B_E666, 32'h432C_CCCC, 32'h432D_B333, 32'h432E_9999, 32'h432F_8000, 32'h4330_6666, 32'h4331_4CCC, 32'h4332_3333, 32'h4332_3333	// 171-179.1
		};

/*		{	32'h0000_0000, 32'h3F80_0000, 32'h4000_0000, 32'h4040_0000, 32'h4080_0000, 32'h40A0_0000, 32'h40C0_0000, 32'h40E0_0000, 32'h4100_0000, 32'h4110_0000,	// 0-9
			32'h4120_0000, 32'h4130_0000, 32'h4140_0000, 32'h4150_0000, 32'h4160_0000, 32'h4170_0000, 32'h4180_0000, 32'h4188_0000, 32'h4190_0000, 32'h4198_0000,	// 10-19
			32'h41A0_0000, 32'h41A8_0000, 32'h41B0_0000, 32'h41B8_0000, 32'h41C0_0000, 32'h41C8_0000, 32'h41D0_0000, 32'h41D8_0000, 32'h41E0_0000, 32'h41E8_0000,	// 20-29
			32'h41F0_0000, 32'h41F8_0000, 32'h4200_0000, 32'h4204_0000, 32'h4208_0000, 32'h420C_0000, 32'h4210_0000, 32'h4214_0000, 32'h4218_0000, 32'h421C_0000,	// 30-39
			32'h4220_0000, 32'h4224_0000, 32'h4228_0000, 32'h422C_0000, 32'h4230_0000, 32'h4234_0000, 32'h4238_0000, 32'h423C_0000, 32'h4240_0000, 32'h4244_0000,	// 40-49
			32'h4248_0000, 32'h424C_0000, 32'h4250_0000, 32'h4254_0000, 32'h4258_0000, 32'h425C_0000, 32'h4260_0000, 32'h4264_0000, 32'h4268_0000, 32'h426C_0000,	// 50-59
			32'h4270_0000, 32'h4274_0000, 32'h4278_0000, 32'h427C_0000, 32'h4280_0000, 32'h4282_0000, 32'h4284_0000, 32'h4286_0000, 32'h4288_0000, 32'h428A_0000,	// 60-69
			32'h428C_0000, 32'h428E_0000, 32'h4290_0000, 32'h4292_0000, 32'h4294_0000, 32'h4296_0000, 32'h4298_0000, 32'h429A_0000, 32'h429C_0000, 32'h429E_0000,	// 70-79
			32'h42A0_0000, 32'h42A2_0000, 32'h42A4_0000, 32'h42A6_0000, 32'h42A8_0000, 32'h42AA_0000, 32'h42AC_0000, 32'h42AE_0000, 32'h42B0_0000, 32'h42B2_0000,	// 80-89
			32'h42B4_0000, 32'h42B6_0000, 32'h42B8_0000, 32'h42BA_0000, 32'h42BC_0000, 32'h42BE_0000, 32'h42C0_0000, 32'h42C2_0000, 32'h42C4_0000, 32'h42C6_0000, 	// 90-99
			32'h42C8_0000, 32'h42CA_0000, 32'h42CC_0000, 32'h42CE_0000, 32'h42D0_0000, 32'h42D2_0000, 32'h42D4_0000, 32'h42D6_0000, 32'h42D8_0000, 32'h42DA_0000, 	// 100-109
			32'h42DC_0000, 32'h42DE_0000, 32'h42E0_0000, 32'h42E2_0000, 32'h42E4_0000, 32'h42E6_0000, 32'h42E8_0000, 32'h42EA_0000, 32'h42EC_0000, 32'h42EE_0000, 	// 110-119
			32'h42F0_0000, 32'h42F2_0000, 32'h42F4_0000, 32'h42F6_0000, 32'h42F8_0000, 32'h42FA_0000, 32'h42FC_0000, 32'h42FE_0000, 32'h4300_0000, 32'h4301_0000, 	// 120-129
			32'h4302_0000, 32'h4303_0000, 32'h4304_0000, 32'h4305_0000, 32'h4306_0000, 32'h4307_0000, 32'h4308_0000, 32'h4309_0000, 32'h430A_0000, 32'h430B_0000, 	// 130-139
			32'h430C_0000, 32'h430D_0000, 32'h430E_0000, 32'h430F_0000, 32'h4310_0000, 32'h4311_0000, 32'h4312_0000, 32'h4313_0000, 32'h4314_0000, 32'h4315_0000, 	// 140-149
			32'h4316_0000, 32'h4317_0000, 32'h4318_0000, 32'h4319_0000, 32'h431A_0000, 32'h431B_0000, 32'h431C_0000, 32'h431D_0000, 32'h431E_0000, 32'h431F_0000, 	// 150-159
			32'h4320_0000, 32'h4321_0000, 32'h4322_0000, 32'h4323_0000, 32'h4324_0000, 32'h4325_0000, 32'h4326_0000, 32'h4327_0000, 32'h4328_0000, 32'h4329_0000, 	// 160-169
			32'h432A_0000, 32'h432B_0000, 32'h432C_0000, 32'h432D_0000, 32'h432E_0000, 32'h432F_0000, 32'h4330_0000, 32'h4331_0000, 32'h4332_0000, 32'h4333_0000	// 170-179
		};
*/

function bit [31:0] sumf;
	input bit [31:0] A, B;
	begin
		if (A == 32'h0000_0000)
			sumf = B;
		else if (B == 32'h0000_0000)
			sumf = A;
		else begin

			sumf[31] = 1'b0;

			if (A[30:23] >= B[30:23]) begin
				sumf[30:23] = B[30:23];
				sumf[22:0] = A[22:0] + (B[22:0] >> (A[30:23] - B[30:23]));
			end
			else begin
				sumf[30:23] = A[30:23];
				sumf[22:0] = B[22:0] + (A[22:0] >> (B[30:23] - A[30:23]));
			end
		end
	end
endfunction
