//--------------------------------------------------------------------------------
//                                                          ������ "���������",���
//                                                          http://www.navigat.ru/
//������    :  
//�����     : CSA
//E-mail    : 
//����      : 
//��������  : ������������ ���� ��� ������ arinc708tx
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
// ����������� ���� ������ arinc708tx 
// ���� �������� ����� 32-� ������ ��������� � ��������� ���������� 
//-------------------------------------------------------------------------------------------------
//
//  �����|  ��� �������� | ��� |  ��������  
//
//  0x00    ID             R      ������� �������������� ���������� ������ � �������  
//  0x01    DATA           R      ��� ������ �� ������� ������ ���������� ������ �� FIFO 
//                                ��������� 32-�������� ����� Arinc 708
//  0x02    NBUF           R      ������� ���������� ���� � FIFO �����������
//  0x03    WBUF           R      ������ FIFO ������   
//  0x04    CTRL           R/W    ������� �������/����������
//  0x05    CSET           W      ������� ����� ��������� � '1' ����� �������� CTRL
//                                ��� ������ ����� �� ������� ������ ������ �� ���� � 
//                                �������� CTRL ��������������� � '1' ,������� �������
//                                ������������� '1' � �����
//                                ��� ������ �� ������� ������ ������������ 'deadbeef'  
//  0x06    CCLR           W      ������� ����� ������ � '0' ����� �������� CTRL
//                                ��� ������ ����� �� ������� ������ ������ �� ���� � 
//                                �������� CTRL ������������ � '0' ,������� �������
//                                ������������� '1' � ����� 
//                                ��� ������ �� ������� ������ ������������ '0xdeadbeef' 
//
//-------------------------------------------------------------------------------------------------
// ������� �������� ��������� 
//-------------------------------------------------------------------------------------------------
// ID:
//      31                              16 15                                 0
//    +-----------------------------------+-----------------------------------+
//    |               ---                 | ������������� ���������� ������   |
//    +-----------------------------------+-----------------------------------+
//    MSB                                                                    LSB
//
// DATA:  ������ ����� Arinc 708, ������������� � FIFO
//    
//      31                              16 15                                 0
//    +-----------------------------------+-----------------------------------+
//    | 							1600 / 32 = 50						      |
//    +-----------------------------------+-----------------------------------+
//    MSB                                                                    LSB
//
//    ���� ������� Arinc708 ���������� 1600 ���. ���� ����������� �� 50 ����
//    �� 32 ������� ������. ����� �������������� � fifo ������
//    ����������� �������� ���� � ���������� ������ -> 0,1,2,3,..,48,49
//    * ��� ������������ ���������� ������ FIFO ������ ��������� ����������� � DATA �     
//     FIFO �� ������������, �� ��������������� ��� ������������ TXF_IF
//    
// CTRL:
//
//        15       14       13       12       11       10       9        8
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//    |TXF_IFD |TXF_IFC |TXF_IFB |TXF_IFA | TXE_FD | TXE_FC | TXE_FB | TXE_FA | ���
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//    |    R   |    R   |    R   |    R   |    R   |    R   |    R   |    R   | ���
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//    |    0   |    0   |    0   |    0   |    0   |   0    |    0   |    0   | ���.����
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//
//        7         6        5        4        3        2        1        0
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//    |  RST   |   --   |   --   |   --   |   --   |   --   |   --   |  ENA   | ���
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//    |  W`1   |   --   |   --   |   --   |   --   |   --   |   --   |   R/W  | ���
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//    |   --   |   --   |   --   |   --   |   --   |   --   |   --   |    0   | ���.����
//    +--------+--------+--------+--------+--------+--------+--------+--------+
//
//    ���: R - ������ �� ������ W - ������ �� ������ R/W - ������ � ������
//         W`1 - ������ ������ ���. 1    
//
//    ENA   -   ���������� ������. ��� ������ ���.1 � ENA ����������� ����� ������

//
//    TXE_FA -  ���� ��������� fifo. ���� ������ ���� ���� ����������, �� �����
//    TXE_FB    ����������� ������ ����� Arinc708
//    TXE_FC
//    TXE_FD
//
//    TXF_IFA - ����  TXF_IF ��������������� � '1' ����� ����� FIFO �������� � ��� ����
//    TXF_IFB   ���������� �������� ������ �� ������ DATA. 
//    TXF_IFC   ���������� ������������ � 0 ��� ������ '1'  �� ������ �� ������� CTRL,CSET,CCLR. 
//    TXF_IFD

    localparam ID      = 0;
    localparam DATA    = 1;
	localparam NBUF    = 2;
	localparam WBUF    = 3;
	localparam CTRL    = 4;
    localparam CSET    = 5;
    localparam CCLR    = 6;		
	
	localparam ENA     = 0;
    localparam RST     = 7;
	
    localparam ADDRESS_DEPTH = 10;
    localparam ADDRESS_WIDTH = 4;
	
    localparam DEFAULT_BDR   = 1_000_000;
	localparam DEFAULT_TMRW  = 100;

	`define ARINC708_FIFO_NWORD	50
	