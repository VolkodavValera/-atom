module UART_Controller (clk, rst_n, rxd, data_rx, data_tx, done);

endmodule // VGA_Controller
