`timescale      1ns / 1ns
`define SYS_CLK 50_000_000

module arinc2vga_tb ();

/*----------------------------------------------------------------------------------*/
/*									Parameters										*/
/*----------------------------------------------------------------------------------*/    
localparam time SYS_CLK_PERIOD = 1_000_000_000.0 / `SYS_CLK;  // (1S-ns / F mhz = P) 

/*----------------------------------------------------------------------------------*/
/*								    Variables										*/
/*----------------------------------------------------------------------------------*/


/*----------------------------------------------------------------------------------*/
/*								Initial blocks										*/
/*----------------------------------------------------------------------------------*/


/*----------------------------------------------------------------------------------*/
/*									Modules											*/
/*----------------------------------------------------------------------------------*/


endmodule